// Generator : SpinalHDL v1.7.3    git head : aeaeece704fe43c766e0d36a93f2ecbb8a9f2003
// Component : dlm_1t2n1c8p
// Git hash  : 69a5423e1bb5ec40bd32371f8e4d623edb0cc7aa

`timescale 1ns/1ps

module dlm_1t2n1c8p (
  input               axi_ctrl_awvalid,
  output              axi_ctrl_awready,
  input      [63:0]   axi_ctrl_awaddr,
  input      [2:0]    axi_ctrl_awprot,
  input               axi_ctrl_wvalid,
  output              axi_ctrl_wready,
  input      [63:0]   axi_ctrl_wdata,
  input      [7:0]    axi_ctrl_wstrb,
  output              axi_ctrl_bvalid,
  input               axi_ctrl_bready,
  output     [1:0]    axi_ctrl_bresp,
  input               axi_ctrl_arvalid,
  output reg          axi_ctrl_arready,
  input      [63:0]   axi_ctrl_araddr,
  input      [2:0]    axi_ctrl_arprot,
  output              axi_ctrl_rvalid,
  input               axi_ctrl_rready,
  output     [63:0]   axi_ctrl_rdata,
  output     [1:0]    axi_ctrl_rresp,
  output              hostd_bpss_rd_req_valid,
  input               hostd_bpss_rd_req_ready,
  output     [95:0]   hostd_bpss_rd_req_data,
  output              hostd_bpss_wr_req_valid,
  input               hostd_bpss_wr_req_ready,
  output     [95:0]   hostd_bpss_wr_req_data,
  input               hostd_bpss_rd_done_valid,
  output              hostd_bpss_rd_done_ready,
  input      [5:0]    hostd_bpss_rd_done_data,
  input               hostd_bpss_wr_done_valid,
  output              hostd_bpss_wr_done_ready,
  input      [5:0]    hostd_bpss_wr_done_data,
  input               hostd_axis_host_sink_tvalid,
  output              hostd_axis_host_sink_tready,
  input      [511:0]  hostd_axis_host_sink_tdata,
  input      [3:0]    hostd_axis_host_sink_tdest,
  input      [63:0]   hostd_axis_host_sink_tkeep,
  input               hostd_axis_host_sink_tlast,
  output              hostd_axis_host_src_tvalid,
  input               hostd_axis_host_src_tready,
  output     [511:0]  hostd_axis_host_src_tdata,
  output     [3:0]    hostd_axis_host_src_tdest,
  output     [63:0]   hostd_axis_host_src_tkeep,
  output              hostd_axis_host_src_tlast,
  output              axi_mem_0_awvalid,
  input               axi_mem_0_awready,
  output     [63:0]   axi_mem_0_awaddr,
  output     [5:0]    axi_mem_0_awid,
  output     [7:0]    axi_mem_0_awlen,
  output     [2:0]    axi_mem_0_awsize,
  output     [1:0]    axi_mem_0_awburst,
  output              axi_mem_0_wvalid,
  input               axi_mem_0_wready,
  output     [511:0]  axi_mem_0_wdata,
  output     [63:0]   axi_mem_0_wstrb,
  output              axi_mem_0_wlast,
  input               axi_mem_0_bvalid,
  output              axi_mem_0_bready,
  input      [5:0]    axi_mem_0_bid,
  input      [1:0]    axi_mem_0_bresp,
  output              axi_mem_0_arvalid,
  input               axi_mem_0_arready,
  output     [63:0]   axi_mem_0_araddr,
  output     [5:0]    axi_mem_0_arid,
  output     [7:0]    axi_mem_0_arlen,
  output     [2:0]    axi_mem_0_arsize,
  output     [1:0]    axi_mem_0_arburst,
  input               axi_mem_0_rvalid,
  output              axi_mem_0_rready,
  input      [511:0]  axi_mem_0_rdata,
  input      [5:0]    axi_mem_0_rid,
  input      [1:0]    axi_mem_0_rresp,
  input               axi_mem_0_rlast,
  output              axi_mem_1_awvalid,
  input               axi_mem_1_awready,
  output     [63:0]   axi_mem_1_awaddr,
  output     [5:0]    axi_mem_1_awid,
  output     [7:0]    axi_mem_1_awlen,
  output     [2:0]    axi_mem_1_awsize,
  output     [1:0]    axi_mem_1_awburst,
  output              axi_mem_1_wvalid,
  input               axi_mem_1_wready,
  output     [511:0]  axi_mem_1_wdata,
  output     [63:0]   axi_mem_1_wstrb,
  output              axi_mem_1_wlast,
  input               axi_mem_1_bvalid,
  output              axi_mem_1_bready,
  input      [5:0]    axi_mem_1_bid,
  input      [1:0]    axi_mem_1_bresp,
  output              axi_mem_1_arvalid,
  input               axi_mem_1_arready,
  output     [63:0]   axi_mem_1_araddr,
  output     [5:0]    axi_mem_1_arid,
  output     [7:0]    axi_mem_1_arlen,
  output     [2:0]    axi_mem_1_arsize,
  output     [1:0]    axi_mem_1_arburst,
  input               axi_mem_1_rvalid,
  output              axi_mem_1_rready,
  input      [511:0]  axi_mem_1_rdata,
  input      [5:0]    axi_mem_1_rid,
  input      [1:0]    axi_mem_1_rresp,
  input               axi_mem_1_rlast,
  output              axi_mem_2_awvalid,
  input               axi_mem_2_awready,
  output     [63:0]   axi_mem_2_awaddr,
  output     [5:0]    axi_mem_2_awid,
  output     [7:0]    axi_mem_2_awlen,
  output     [2:0]    axi_mem_2_awsize,
  output     [1:0]    axi_mem_2_awburst,
  output              axi_mem_2_wvalid,
  input               axi_mem_2_wready,
  output     [511:0]  axi_mem_2_wdata,
  output     [63:0]   axi_mem_2_wstrb,
  output              axi_mem_2_wlast,
  input               axi_mem_2_bvalid,
  output              axi_mem_2_bready,
  input      [5:0]    axi_mem_2_bid,
  input      [1:0]    axi_mem_2_bresp,
  output              axi_mem_2_arvalid,
  input               axi_mem_2_arready,
  output     [63:0]   axi_mem_2_araddr,
  output     [5:0]    axi_mem_2_arid,
  output     [7:0]    axi_mem_2_arlen,
  output     [2:0]    axi_mem_2_arsize,
  output     [1:0]    axi_mem_2_arburst,
  input               axi_mem_2_rvalid,
  output              axi_mem_2_rready,
  input      [511:0]  axi_mem_2_rdata,
  input      [5:0]    axi_mem_2_rid,
  input      [1:0]    axi_mem_2_rresp,
  input               axi_mem_2_rlast,
  output              axi_mem_3_awvalid,
  input               axi_mem_3_awready,
  output     [63:0]   axi_mem_3_awaddr,
  output     [5:0]    axi_mem_3_awid,
  output     [7:0]    axi_mem_3_awlen,
  output     [2:0]    axi_mem_3_awsize,
  output     [1:0]    axi_mem_3_awburst,
  output              axi_mem_3_wvalid,
  input               axi_mem_3_wready,
  output     [511:0]  axi_mem_3_wdata,
  output     [63:0]   axi_mem_3_wstrb,
  output              axi_mem_3_wlast,
  input               axi_mem_3_bvalid,
  output              axi_mem_3_bready,
  input      [5:0]    axi_mem_3_bid,
  input      [1:0]    axi_mem_3_bresp,
  output              axi_mem_3_arvalid,
  input               axi_mem_3_arready,
  output     [63:0]   axi_mem_3_araddr,
  output     [5:0]    axi_mem_3_arid,
  output     [7:0]    axi_mem_3_arlen,
  output     [2:0]    axi_mem_3_arsize,
  output     [1:0]    axi_mem_3_arburst,
  input               axi_mem_3_rvalid,
  output              axi_mem_3_rready,
  input      [511:0]  axi_mem_3_rdata,
  input      [5:0]    axi_mem_3_rid,
  input      [1:0]    axi_mem_3_rresp,
  input               axi_mem_3_rlast,
  input               rdma_0_rd_req_valid,
  output              rdma_0_rd_req_ready,
  input      [95:0]   rdma_0_rd_req_data,
  input               rdma_0_wr_req_valid,
  output              rdma_0_wr_req_ready,
  input      [95:0]   rdma_0_wr_req_data,
  output              rdma_0_sq_valid,
  input               rdma_0_sq_ready,
  output     [543:0]  rdma_0_sq_data,
  input               rdma_0_ack_valid,
  output              rdma_0_ack_ready,
  input      [42:0]   rdma_0_ack_data,
  input               rdma_0_axis_sink_tvalid,
  output              rdma_0_axis_sink_tready,
  input      [511:0]  rdma_0_axis_sink_tdata,
  input      [63:0]   rdma_0_axis_sink_tkeep,
  input               rdma_0_axis_sink_tlast,
  output              rdma_0_axis_src_tvalid,
  input               rdma_0_axis_src_tready,
  output     [511:0]  rdma_0_axis_src_tdata,
  output     [63:0]   rdma_0_axis_src_tkeep,
  output              rdma_0_axis_src_tlast,
  input               resetn,
  input               clk
);

  wire       [63:0]   hbmHost_io_cntDone;
  wire                hbmHost_io_hostd_bpss_rd_req_valid;
  wire       [95:0]   hbmHost_io_hostd_bpss_rd_req_payload_data;
  wire                hbmHost_io_hostd_bpss_wr_req_valid;
  wire       [95:0]   hbmHost_io_hostd_bpss_wr_req_payload_data;
  wire                hbmHost_io_hostd_bpss_rd_done_ready;
  wire                hbmHost_io_hostd_bpss_wr_done_ready;
  wire                hbmHost_io_hostd_axis_host_sink_ready;
  wire                hbmHost_io_hostd_axis_host_src_valid;
  wire       [511:0]  hbmHost_io_hostd_axis_host_src_payload_tdata;
  wire       [3:0]    hbmHost_io_hostd_axis_host_src_payload_tdest;
  wire       [63:0]   hbmHost_io_hostd_axis_host_src_payload_tkeep;
  wire                hbmHost_io_hostd_axis_host_src_payload_tlast;
  wire                hbmHost_io_axi_cmem_ar_valid;
  wire       [63:0]   hbmHost_io_axi_cmem_ar_payload_addr;
  wire       [5:0]    hbmHost_io_axi_cmem_ar_payload_id;
  wire       [7:0]    hbmHost_io_axi_cmem_ar_payload_len;
  wire       [2:0]    hbmHost_io_axi_cmem_ar_payload_size;
  wire       [1:0]    hbmHost_io_axi_cmem_ar_payload_burst;
  wire                hbmHost_io_axi_cmem_aw_valid;
  wire       [63:0]   hbmHost_io_axi_cmem_aw_payload_addr;
  wire       [5:0]    hbmHost_io_axi_cmem_aw_payload_id;
  wire       [7:0]    hbmHost_io_axi_cmem_aw_payload_len;
  wire       [2:0]    hbmHost_io_axi_cmem_aw_payload_size;
  wire       [1:0]    hbmHost_io_axi_cmem_aw_payload_burst;
  wire                hbmHost_io_axi_cmem_w_valid;
  wire       [511:0]  hbmHost_io_axi_cmem_w_payload_data;
  wire       [63:0]   hbmHost_io_axi_cmem_w_payload_strb;
  wire                hbmHost_io_axi_cmem_w_payload_last;
  wire                hbmHost_io_axi_cmem_r_ready;
  wire                hbmHost_io_axi_cmem_b_ready;
  wire                txnEng_io_node_axi_0_ar_valid;
  wire       [63:0]   txnEng_io_node_axi_0_ar_payload_addr;
  wire       [5:0]    txnEng_io_node_axi_0_ar_payload_id;
  wire       [7:0]    txnEng_io_node_axi_0_ar_payload_len;
  wire       [2:0]    txnEng_io_node_axi_0_ar_payload_size;
  wire       [1:0]    txnEng_io_node_axi_0_ar_payload_burst;
  wire                txnEng_io_node_axi_0_aw_valid;
  wire       [63:0]   txnEng_io_node_axi_0_aw_payload_addr;
  wire       [5:0]    txnEng_io_node_axi_0_aw_payload_id;
  wire       [7:0]    txnEng_io_node_axi_0_aw_payload_len;
  wire       [2:0]    txnEng_io_node_axi_0_aw_payload_size;
  wire       [1:0]    txnEng_io_node_axi_0_aw_payload_burst;
  wire                txnEng_io_node_axi_0_w_valid;
  wire       [511:0]  txnEng_io_node_axi_0_w_payload_data;
  wire       [63:0]   txnEng_io_node_axi_0_w_payload_strb;
  wire                txnEng_io_node_axi_0_w_payload_last;
  wire                txnEng_io_node_axi_0_r_ready;
  wire                txnEng_io_node_axi_0_b_ready;
  wire                txnEng_io_node_axi_1_ar_valid;
  wire       [63:0]   txnEng_io_node_axi_1_ar_payload_addr;
  wire       [5:0]    txnEng_io_node_axi_1_ar_payload_id;
  wire       [7:0]    txnEng_io_node_axi_1_ar_payload_len;
  wire       [2:0]    txnEng_io_node_axi_1_ar_payload_size;
  wire       [1:0]    txnEng_io_node_axi_1_ar_payload_burst;
  wire                txnEng_io_node_axi_1_aw_valid;
  wire       [63:0]   txnEng_io_node_axi_1_aw_payload_addr;
  wire       [5:0]    txnEng_io_node_axi_1_aw_payload_id;
  wire       [7:0]    txnEng_io_node_axi_1_aw_payload_len;
  wire       [2:0]    txnEng_io_node_axi_1_aw_payload_size;
  wire       [1:0]    txnEng_io_node_axi_1_aw_payload_burst;
  wire                txnEng_io_node_axi_1_w_valid;
  wire       [511:0]  txnEng_io_node_axi_1_w_payload_data;
  wire       [63:0]   txnEng_io_node_axi_1_w_payload_strb;
  wire                txnEng_io_node_axi_1_w_payload_last;
  wire                txnEng_io_node_axi_1_r_ready;
  wire                txnEng_io_node_axi_1_b_ready;
  wire                txnEng_io_node_cmdAxi_0_ar_valid;
  wire       [63:0]   txnEng_io_node_cmdAxi_0_ar_payload_addr;
  wire       [5:0]    txnEng_io_node_cmdAxi_0_ar_payload_id;
  wire       [7:0]    txnEng_io_node_cmdAxi_0_ar_payload_len;
  wire       [2:0]    txnEng_io_node_cmdAxi_0_ar_payload_size;
  wire       [1:0]    txnEng_io_node_cmdAxi_0_ar_payload_burst;
  wire                txnEng_io_node_cmdAxi_0_aw_valid;
  wire       [63:0]   txnEng_io_node_cmdAxi_0_aw_payload_addr;
  wire       [5:0]    txnEng_io_node_cmdAxi_0_aw_payload_id;
  wire       [7:0]    txnEng_io_node_cmdAxi_0_aw_payload_len;
  wire       [2:0]    txnEng_io_node_cmdAxi_0_aw_payload_size;
  wire       [1:0]    txnEng_io_node_cmdAxi_0_aw_payload_burst;
  wire                txnEng_io_node_cmdAxi_0_w_valid;
  wire       [511:0]  txnEng_io_node_cmdAxi_0_w_payload_data;
  wire       [63:0]   txnEng_io_node_cmdAxi_0_w_payload_strb;
  wire                txnEng_io_node_cmdAxi_0_w_payload_last;
  wire                txnEng_io_node_cmdAxi_0_r_ready;
  wire                txnEng_io_node_cmdAxi_0_b_ready;
  wire                txnEng_io_node_done_0;
  wire       [31:0]   txnEng_io_node_cntTxnCmt_0;
  wire       [31:0]   txnEng_io_node_cntTxnAbt_0;
  wire       [31:0]   txnEng_io_node_cntTxnLd_0;
  wire       [31:0]   txnEng_io_node_cntLockLoc_0;
  wire       [31:0]   txnEng_io_node_cntLockRmt_0;
  wire       [31:0]   txnEng_io_node_cntLockDenyLoc_0;
  wire       [31:0]   txnEng_io_node_cntLockDenyRmt_0;
  wire       [31:0]   txnEng_io_node_cntClk_0;
  wire                txnEng_io_rdma_rd_req_ready;
  wire                txnEng_io_rdma_wr_req_ready;
  wire                txnEng_io_rdma_sq_valid;
  wire       [543:0]  txnEng_io_rdma_sq_payload_data;
  wire                txnEng_io_rdma_ack_ready;
  wire                txnEng_io_rdma_axis_sink_ready;
  wire                txnEng_io_rdma_axis_src_valid;
  wire       [511:0]  txnEng_io_rdma_axis_src_payload_tdata;
  wire       [63:0]   txnEng_io_rdma_axis_src_payload_tkeep;
  wire                txnEng_io_rdma_axis_src_payload_tlast;
  wire       [31:0]   txnEng_io_cntRDMASent;
  wire       [31:0]   txnEng_io_cntRDMARecv;
  wire                ctrlR_readHaltRequest;
  wire                ctrlR_writeHaltRequest;
  wire                ctrlR_writeJoinEvent_valid;
  wire                ctrlR_writeJoinEvent_ready;
  wire                ctrlR_writeJoinEvent_fire;
  wire       [1:0]    ctrlR_writeRsp_resp;
  wire                ctrlR_writeJoinEvent_translated_valid;
  wire                ctrlR_writeJoinEvent_translated_ready;
  wire       [1:0]    ctrlR_writeJoinEvent_translated_payload_resp;
  wire                _zz_axi_ctrl_bvalid;
  reg                 _zz_ctrlR_writeJoinEvent_translated_ready;
  wire                _zz_axi_ctrl_bvalid_1;
  reg                 _zz_axi_ctrl_bvalid_2;
  reg        [1:0]    _zz_axi_ctrl_bresp;
  wire                when_Stream_l368;
  wire                ctrlR_readDataStage_valid;
  wire                ctrlR_readDataStage_ready;
  wire       [63:0]   ctrlR_readDataStage_payload_addr;
  wire       [2:0]    ctrlR_readDataStage_payload_prot;
  reg                 axi_ctrl_ar_rValid;
  reg        [63:0]   axi_ctrl_ar_rData_addr;
  reg        [2:0]    axi_ctrl_ar_rData_prot;
  wire                when_Stream_l368_1;
  reg        [63:0]   ctrlR_readRsp_data;
  wire       [1:0]    ctrlR_readRsp_resp;
  wire                _zz_axi_ctrl_rvalid;
  wire       [63:0]   ctrlR_readAddressMasked;
  wire       [63:0]   ctrlR_writeAddressMasked;
  wire                ctrlR_writeOccur;
  wire                ctrlR_readOccur;
  reg        [1:0]    _zz_ctrlR_readRsp_data;
  wire                when_Types_l264;
  reg        [63:0]   _zz_ctrlR_readRsp_data_1;
  reg        [63:0]   _zz_ctrlR_readRsp_data_2;
  reg        [15:0]   _zz_ctrlR_readRsp_data_3;
  reg        [63:0]   _zz_ctrlR_readRsp_data_4;
  reg        [5:0]    _zz_ctrlR_readRsp_data_5;
  reg                 _zz_ctrlR_readRsp_data_6;
  reg        [31:0]   _zz_ctrlR_readRsp_data_7;
  reg        [9:0]    _zz_ctrlR_readRsp_data_8;
  reg        [3:0]    _zz_ctrlR_readRsp_data_9;
  reg                 _zz_ctrlR_readRsp_data_10;
  reg        [31:0]   _zz_ctrlR_readRsp_data_11;
  reg        [9:0]    _zz_ctrlR_readRsp_data_12;
  reg        [3:0]    _zz_ctrlR_readRsp_data_13;
  reg                 when_Types_l284;
  reg        [0:0]    _zz_ctrlR_readRsp_data_14;
  reg        [31:0]   _zz_ctrlR_readRsp_data_15;
  reg        [31:0]   _zz_ctrlR_readRsp_data_16;
  wire                when_BusSlaveFactory_l962;
  wire                when_BusSlaveFactory_l962_1;
  wire                when_BusSlaveFactory_l962_2;
  wire                when_BusSlaveFactory_l962_3;
  wire                when_BusSlaveFactory_l962_4;
  wire                when_BusSlaveFactory_l962_5;
  wire                when_BusSlaveFactory_l962_6;
  wire                when_BusSlaveFactory_l962_7;
  wire                when_BusSlaveFactory_l962_8;
  wire                when_BusSlaveFactory_l962_9;
  wire                when_BusSlaveFactory_l962_10;
  wire                when_BusSlaveFactory_l962_11;
  wire                when_BusSlaveFactory_l962_12;
  wire                when_BusSlaveFactory_l962_13;
  wire                when_BusSlaveFactory_l962_14;
  wire                when_BusSlaveFactory_l962_15;
  wire                when_BusSlaveFactory_l962_16;
  wire                when_BusSlaveFactory_l962_17;
  wire                when_BusSlaveFactory_l962_18;
  wire                when_BusSlaveFactory_l962_19;
  wire                when_BusSlaveFactory_l962_20;
  wire                when_BusSlaveFactory_l962_21;
  wire                when_BusSlaveFactory_l962_22;
  wire                when_BusSlaveFactory_l962_23;
  wire                when_BusSlaveFactory_l962_24;
  wire                when_BusSlaveFactory_l962_25;
  wire                when_BusSlaveFactory_l962_26;
  wire                when_BusSlaveFactory_l962_27;
  wire                when_BusSlaveFactory_l962_28;
  wire                when_BusSlaveFactory_l962_29;
  wire                when_BusSlaveFactory_l962_30;
  wire                when_BusSlaveFactory_l962_31;
  wire                when_BusSlaveFactory_l962_32;
  wire                when_BusSlaveFactory_l962_33;
  wire                when_BusSlaveFactory_l962_34;
  wire                when_BusSlaveFactory_l962_35;
  wire                when_BusSlaveFactory_l962_36;
  wire                when_BusSlaveFactory_l962_37;
  wire                when_BusSlaveFactory_l962_38;
  wire                when_BusSlaveFactory_l962_39;
  wire                when_BusSlaveFactory_l962_40;
  wire                when_BusSlaveFactory_l962_41;
  wire                when_BusSlaveFactory_l962_42;
  wire                when_BusSlaveFactory_l962_43;
  wire                when_BusSlaveFactory_l962_44;
  wire                when_BusSlaveFactory_l962_45;
  wire                when_BusSlaveFactory_l962_46;
  wire                when_BusSlaveFactory_l962_47;
  wire                when_BusSlaveFactory_l962_48;
  wire                when_BusSlaveFactory_l962_49;
  wire                when_BusSlaveFactory_l962_50;
  wire                when_BusSlaveFactory_l962_51;
  wire                when_BusSlaveFactory_l962_52;
  wire                when_BusSlaveFactory_l962_53;
  wire                when_BusSlaveFactory_l962_54;
  wire                when_BusSlaveFactory_l962_55;

  CMemHost hbmHost (
    .io_mode                               (_zz_ctrlR_readRsp_data[1:0]                        ), //i
    .io_hostAddr                           (_zz_ctrlR_readRsp_data_1[63:0]                     ), //i
    .io_cmemAddr                           (_zz_ctrlR_readRsp_data_2[63:0]                     ), //i
    .io_len                                (_zz_ctrlR_readRsp_data_3[15:0]                     ), //i
    .io_cnt                                (_zz_ctrlR_readRsp_data_4[63:0]                     ), //i
    .io_pid                                (_zz_ctrlR_readRsp_data_5[5:0]                      ), //i
    .io_cntDone                            (hbmHost_io_cntDone[63:0]                           ), //o
    .io_hostd_bpss_rd_req_valid            (hbmHost_io_hostd_bpss_rd_req_valid                 ), //o
    .io_hostd_bpss_rd_req_ready            (hostd_bpss_rd_req_ready                            ), //i
    .io_hostd_bpss_rd_req_payload_data     (hbmHost_io_hostd_bpss_rd_req_payload_data[95:0]    ), //o
    .io_hostd_bpss_wr_req_valid            (hbmHost_io_hostd_bpss_wr_req_valid                 ), //o
    .io_hostd_bpss_wr_req_ready            (hostd_bpss_wr_req_ready                            ), //i
    .io_hostd_bpss_wr_req_payload_data     (hbmHost_io_hostd_bpss_wr_req_payload_data[95:0]    ), //o
    .io_hostd_bpss_rd_done_valid           (hostd_bpss_rd_done_valid                           ), //i
    .io_hostd_bpss_rd_done_ready           (hbmHost_io_hostd_bpss_rd_done_ready                ), //o
    .io_hostd_bpss_rd_done_payload_data    (hostd_bpss_rd_done_data[5:0]                       ), //i
    .io_hostd_bpss_wr_done_valid           (hostd_bpss_wr_done_valid                           ), //i
    .io_hostd_bpss_wr_done_ready           (hbmHost_io_hostd_bpss_wr_done_ready                ), //o
    .io_hostd_bpss_wr_done_payload_data    (hostd_bpss_wr_done_data[5:0]                       ), //i
    .io_hostd_axis_host_sink_valid         (hostd_axis_host_sink_tvalid                        ), //i
    .io_hostd_axis_host_sink_ready         (hbmHost_io_hostd_axis_host_sink_ready              ), //o
    .io_hostd_axis_host_sink_payload_tdata (hostd_axis_host_sink_tdata[511:0]                  ), //i
    .io_hostd_axis_host_sink_payload_tdest (hostd_axis_host_sink_tdest[3:0]                    ), //i
    .io_hostd_axis_host_sink_payload_tkeep (hostd_axis_host_sink_tkeep[63:0]                   ), //i
    .io_hostd_axis_host_sink_payload_tlast (hostd_axis_host_sink_tlast                         ), //i
    .io_hostd_axis_host_src_valid          (hbmHost_io_hostd_axis_host_src_valid               ), //o
    .io_hostd_axis_host_src_ready          (hostd_axis_host_src_tready                         ), //i
    .io_hostd_axis_host_src_payload_tdata  (hbmHost_io_hostd_axis_host_src_payload_tdata[511:0]), //o
    .io_hostd_axis_host_src_payload_tdest  (hbmHost_io_hostd_axis_host_src_payload_tdest[3:0]  ), //o
    .io_hostd_axis_host_src_payload_tkeep  (hbmHost_io_hostd_axis_host_src_payload_tkeep[63:0] ), //o
    .io_hostd_axis_host_src_payload_tlast  (hbmHost_io_hostd_axis_host_src_payload_tlast       ), //o
    .io_axi_cmem_aw_valid                  (hbmHost_io_axi_cmem_aw_valid                       ), //o
    .io_axi_cmem_aw_ready                  (axi_mem_0_awready                                  ), //i
    .io_axi_cmem_aw_payload_addr           (hbmHost_io_axi_cmem_aw_payload_addr[63:0]          ), //o
    .io_axi_cmem_aw_payload_id             (hbmHost_io_axi_cmem_aw_payload_id[5:0]             ), //o
    .io_axi_cmem_aw_payload_len            (hbmHost_io_axi_cmem_aw_payload_len[7:0]            ), //o
    .io_axi_cmem_aw_payload_size           (hbmHost_io_axi_cmem_aw_payload_size[2:0]           ), //o
    .io_axi_cmem_aw_payload_burst          (hbmHost_io_axi_cmem_aw_payload_burst[1:0]          ), //o
    .io_axi_cmem_w_valid                   (hbmHost_io_axi_cmem_w_valid                        ), //o
    .io_axi_cmem_w_ready                   (axi_mem_0_wready                                   ), //i
    .io_axi_cmem_w_payload_data            (hbmHost_io_axi_cmem_w_payload_data[511:0]          ), //o
    .io_axi_cmem_w_payload_strb            (hbmHost_io_axi_cmem_w_payload_strb[63:0]           ), //o
    .io_axi_cmem_w_payload_last            (hbmHost_io_axi_cmem_w_payload_last                 ), //o
    .io_axi_cmem_b_valid                   (axi_mem_0_bvalid                                   ), //i
    .io_axi_cmem_b_ready                   (hbmHost_io_axi_cmem_b_ready                        ), //o
    .io_axi_cmem_b_payload_id              (axi_mem_0_bid[5:0]                                 ), //i
    .io_axi_cmem_b_payload_resp            (axi_mem_0_bresp[1:0]                               ), //i
    .io_axi_cmem_ar_valid                  (hbmHost_io_axi_cmem_ar_valid                       ), //o
    .io_axi_cmem_ar_ready                  (axi_mem_0_arready                                  ), //i
    .io_axi_cmem_ar_payload_addr           (hbmHost_io_axi_cmem_ar_payload_addr[63:0]          ), //o
    .io_axi_cmem_ar_payload_id             (hbmHost_io_axi_cmem_ar_payload_id[5:0]             ), //o
    .io_axi_cmem_ar_payload_len            (hbmHost_io_axi_cmem_ar_payload_len[7:0]            ), //o
    .io_axi_cmem_ar_payload_size           (hbmHost_io_axi_cmem_ar_payload_size[2:0]           ), //o
    .io_axi_cmem_ar_payload_burst          (hbmHost_io_axi_cmem_ar_payload_burst[1:0]          ), //o
    .io_axi_cmem_r_valid                   (axi_mem_0_rvalid                                   ), //i
    .io_axi_cmem_r_ready                   (hbmHost_io_axi_cmem_r_ready                        ), //o
    .io_axi_cmem_r_payload_data            (axi_mem_0_rdata[511:0]                             ), //i
    .io_axi_cmem_r_payload_id              (axi_mem_0_rid[5:0]                                 ), //i
    .io_axi_cmem_r_payload_resp            (axi_mem_0_rresp[1:0]                               ), //i
    .io_axi_cmem_r_payload_last            (axi_mem_0_rlast                                    ), //i
    .clk                                   (clk                                                ), //i
    .resetn                                (resetn                                             )  //i
  );
  WrapNodeNet txnEng (
    .io_node_axi_0_aw_valid            (txnEng_io_node_axi_0_aw_valid                ), //o
    .io_node_axi_0_aw_ready            (axi_mem_1_awready                            ), //i
    .io_node_axi_0_aw_payload_addr     (txnEng_io_node_axi_0_aw_payload_addr[63:0]   ), //o
    .io_node_axi_0_aw_payload_id       (txnEng_io_node_axi_0_aw_payload_id[5:0]      ), //o
    .io_node_axi_0_aw_payload_len      (txnEng_io_node_axi_0_aw_payload_len[7:0]     ), //o
    .io_node_axi_0_aw_payload_size     (txnEng_io_node_axi_0_aw_payload_size[2:0]    ), //o
    .io_node_axi_0_aw_payload_burst    (txnEng_io_node_axi_0_aw_payload_burst[1:0]   ), //o
    .io_node_axi_0_w_valid             (txnEng_io_node_axi_0_w_valid                 ), //o
    .io_node_axi_0_w_ready             (axi_mem_1_wready                             ), //i
    .io_node_axi_0_w_payload_data      (txnEng_io_node_axi_0_w_payload_data[511:0]   ), //o
    .io_node_axi_0_w_payload_strb      (txnEng_io_node_axi_0_w_payload_strb[63:0]    ), //o
    .io_node_axi_0_w_payload_last      (txnEng_io_node_axi_0_w_payload_last          ), //o
    .io_node_axi_0_b_valid             (axi_mem_1_bvalid                             ), //i
    .io_node_axi_0_b_ready             (txnEng_io_node_axi_0_b_ready                 ), //o
    .io_node_axi_0_b_payload_id        (axi_mem_1_bid[5:0]                           ), //i
    .io_node_axi_0_b_payload_resp      (axi_mem_1_bresp[1:0]                         ), //i
    .io_node_axi_0_ar_valid            (txnEng_io_node_axi_0_ar_valid                ), //o
    .io_node_axi_0_ar_ready            (axi_mem_1_arready                            ), //i
    .io_node_axi_0_ar_payload_addr     (txnEng_io_node_axi_0_ar_payload_addr[63:0]   ), //o
    .io_node_axi_0_ar_payload_id       (txnEng_io_node_axi_0_ar_payload_id[5:0]      ), //o
    .io_node_axi_0_ar_payload_len      (txnEng_io_node_axi_0_ar_payload_len[7:0]     ), //o
    .io_node_axi_0_ar_payload_size     (txnEng_io_node_axi_0_ar_payload_size[2:0]    ), //o
    .io_node_axi_0_ar_payload_burst    (txnEng_io_node_axi_0_ar_payload_burst[1:0]   ), //o
    .io_node_axi_0_r_valid             (axi_mem_1_rvalid                             ), //i
    .io_node_axi_0_r_ready             (txnEng_io_node_axi_0_r_ready                 ), //o
    .io_node_axi_0_r_payload_data      (axi_mem_1_rdata[511:0]                       ), //i
    .io_node_axi_0_r_payload_id        (axi_mem_1_rid[5:0]                           ), //i
    .io_node_axi_0_r_payload_resp      (axi_mem_1_rresp[1:0]                         ), //i
    .io_node_axi_0_r_payload_last      (axi_mem_1_rlast                              ), //i
    .io_node_axi_1_aw_valid            (txnEng_io_node_axi_1_aw_valid                ), //o
    .io_node_axi_1_aw_ready            (axi_mem_2_awready                            ), //i
    .io_node_axi_1_aw_payload_addr     (txnEng_io_node_axi_1_aw_payload_addr[63:0]   ), //o
    .io_node_axi_1_aw_payload_id       (txnEng_io_node_axi_1_aw_payload_id[5:0]      ), //o
    .io_node_axi_1_aw_payload_len      (txnEng_io_node_axi_1_aw_payload_len[7:0]     ), //o
    .io_node_axi_1_aw_payload_size     (txnEng_io_node_axi_1_aw_payload_size[2:0]    ), //o
    .io_node_axi_1_aw_payload_burst    (txnEng_io_node_axi_1_aw_payload_burst[1:0]   ), //o
    .io_node_axi_1_w_valid             (txnEng_io_node_axi_1_w_valid                 ), //o
    .io_node_axi_1_w_ready             (axi_mem_2_wready                             ), //i
    .io_node_axi_1_w_payload_data      (txnEng_io_node_axi_1_w_payload_data[511:0]   ), //o
    .io_node_axi_1_w_payload_strb      (txnEng_io_node_axi_1_w_payload_strb[63:0]    ), //o
    .io_node_axi_1_w_payload_last      (txnEng_io_node_axi_1_w_payload_last          ), //o
    .io_node_axi_1_b_valid             (axi_mem_2_bvalid                             ), //i
    .io_node_axi_1_b_ready             (txnEng_io_node_axi_1_b_ready                 ), //o
    .io_node_axi_1_b_payload_id        (axi_mem_2_bid[5:0]                           ), //i
    .io_node_axi_1_b_payload_resp      (axi_mem_2_bresp[1:0]                         ), //i
    .io_node_axi_1_ar_valid            (txnEng_io_node_axi_1_ar_valid                ), //o
    .io_node_axi_1_ar_ready            (axi_mem_2_arready                            ), //i
    .io_node_axi_1_ar_payload_addr     (txnEng_io_node_axi_1_ar_payload_addr[63:0]   ), //o
    .io_node_axi_1_ar_payload_id       (txnEng_io_node_axi_1_ar_payload_id[5:0]      ), //o
    .io_node_axi_1_ar_payload_len      (txnEng_io_node_axi_1_ar_payload_len[7:0]     ), //o
    .io_node_axi_1_ar_payload_size     (txnEng_io_node_axi_1_ar_payload_size[2:0]    ), //o
    .io_node_axi_1_ar_payload_burst    (txnEng_io_node_axi_1_ar_payload_burst[1:0]   ), //o
    .io_node_axi_1_r_valid             (axi_mem_2_rvalid                             ), //i
    .io_node_axi_1_r_ready             (txnEng_io_node_axi_1_r_ready                 ), //o
    .io_node_axi_1_r_payload_data      (axi_mem_2_rdata[511:0]                       ), //i
    .io_node_axi_1_r_payload_id        (axi_mem_2_rid[5:0]                           ), //i
    .io_node_axi_1_r_payload_resp      (axi_mem_2_rresp[1:0]                         ), //i
    .io_node_axi_1_r_payload_last      (axi_mem_2_rlast                              ), //i
    .io_node_cmdAxi_0_aw_valid         (txnEng_io_node_cmdAxi_0_aw_valid             ), //o
    .io_node_cmdAxi_0_aw_ready         (axi_mem_3_awready                            ), //i
    .io_node_cmdAxi_0_aw_payload_addr  (txnEng_io_node_cmdAxi_0_aw_payload_addr[63:0]), //o
    .io_node_cmdAxi_0_aw_payload_id    (txnEng_io_node_cmdAxi_0_aw_payload_id[5:0]   ), //o
    .io_node_cmdAxi_0_aw_payload_len   (txnEng_io_node_cmdAxi_0_aw_payload_len[7:0]  ), //o
    .io_node_cmdAxi_0_aw_payload_size  (txnEng_io_node_cmdAxi_0_aw_payload_size[2:0] ), //o
    .io_node_cmdAxi_0_aw_payload_burst (txnEng_io_node_cmdAxi_0_aw_payload_burst[1:0]), //o
    .io_node_cmdAxi_0_w_valid          (txnEng_io_node_cmdAxi_0_w_valid              ), //o
    .io_node_cmdAxi_0_w_ready          (axi_mem_3_wready                             ), //i
    .io_node_cmdAxi_0_w_payload_data   (txnEng_io_node_cmdAxi_0_w_payload_data[511:0]), //o
    .io_node_cmdAxi_0_w_payload_strb   (txnEng_io_node_cmdAxi_0_w_payload_strb[63:0] ), //o
    .io_node_cmdAxi_0_w_payload_last   (txnEng_io_node_cmdAxi_0_w_payload_last       ), //o
    .io_node_cmdAxi_0_b_valid          (axi_mem_3_bvalid                             ), //i
    .io_node_cmdAxi_0_b_ready          (txnEng_io_node_cmdAxi_0_b_ready              ), //o
    .io_node_cmdAxi_0_b_payload_id     (axi_mem_3_bid[5:0]                           ), //i
    .io_node_cmdAxi_0_b_payload_resp   (axi_mem_3_bresp[1:0]                         ), //i
    .io_node_cmdAxi_0_ar_valid         (txnEng_io_node_cmdAxi_0_ar_valid             ), //o
    .io_node_cmdAxi_0_ar_ready         (axi_mem_3_arready                            ), //i
    .io_node_cmdAxi_0_ar_payload_addr  (txnEng_io_node_cmdAxi_0_ar_payload_addr[63:0]), //o
    .io_node_cmdAxi_0_ar_payload_id    (txnEng_io_node_cmdAxi_0_ar_payload_id[5:0]   ), //o
    .io_node_cmdAxi_0_ar_payload_len   (txnEng_io_node_cmdAxi_0_ar_payload_len[7:0]  ), //o
    .io_node_cmdAxi_0_ar_payload_size  (txnEng_io_node_cmdAxi_0_ar_payload_size[2:0] ), //o
    .io_node_cmdAxi_0_ar_payload_burst (txnEng_io_node_cmdAxi_0_ar_payload_burst[1:0]), //o
    .io_node_cmdAxi_0_r_valid          (axi_mem_3_rvalid                             ), //i
    .io_node_cmdAxi_0_r_ready          (txnEng_io_node_cmdAxi_0_r_ready              ), //o
    .io_node_cmdAxi_0_r_payload_data   (axi_mem_3_rdata[511:0]                       ), //i
    .io_node_cmdAxi_0_r_payload_id     (axi_mem_3_rid[5:0]                           ), //i
    .io_node_cmdAxi_0_r_payload_resp   (axi_mem_3_rresp[1:0]                         ), //i
    .io_node_cmdAxi_0_r_payload_last   (axi_mem_3_rlast                              ), //i
    .io_node_nodeId                    (_zz_ctrlR_readRsp_data_14                    ), //i
    .io_node_txnNumTotal               (_zz_ctrlR_readRsp_data_15[31:0]              ), //i
    .io_node_cmdAddrOffs_0             (_zz_ctrlR_readRsp_data_16[31:0]              ), //i
    .io_node_start                     (when_Types_l284                              ), //i
    .io_node_done_0                    (txnEng_io_node_done_0                        ), //o
    .io_node_cntTxnCmt_0               (txnEng_io_node_cntTxnCmt_0[31:0]             ), //o
    .io_node_cntTxnAbt_0               (txnEng_io_node_cntTxnAbt_0[31:0]             ), //o
    .io_node_cntTxnLd_0                (txnEng_io_node_cntTxnLd_0[31:0]              ), //o
    .io_node_cntLockLoc_0              (txnEng_io_node_cntLockLoc_0[31:0]            ), //o
    .io_node_cntLockRmt_0              (txnEng_io_node_cntLockRmt_0[31:0]            ), //o
    .io_node_cntLockDenyLoc_0          (txnEng_io_node_cntLockDenyLoc_0[31:0]        ), //o
    .io_node_cntLockDenyRmt_0          (txnEng_io_node_cntLockDenyRmt_0[31:0]        ), //o
    .io_node_cntClk_0                  (txnEng_io_node_cntClk_0[31:0]                ), //o
    .io_rdma_rd_req_valid              (rdma_0_rd_req_valid                          ), //i
    .io_rdma_rd_req_ready              (txnEng_io_rdma_rd_req_ready                  ), //o
    .io_rdma_rd_req_payload_data       (rdma_0_rd_req_data[95:0]                     ), //i
    .io_rdma_wr_req_valid              (rdma_0_wr_req_valid                          ), //i
    .io_rdma_wr_req_ready              (txnEng_io_rdma_wr_req_ready                  ), //o
    .io_rdma_wr_req_payload_data       (rdma_0_wr_req_data[95:0]                     ), //i
    .io_rdma_sq_valid                  (txnEng_io_rdma_sq_valid                      ), //o
    .io_rdma_sq_ready                  (rdma_0_sq_ready                              ), //i
    .io_rdma_sq_payload_data           (txnEng_io_rdma_sq_payload_data[543:0]        ), //o
    .io_rdma_ack_valid                 (rdma_0_ack_valid                             ), //i
    .io_rdma_ack_ready                 (txnEng_io_rdma_ack_ready                     ), //o
    .io_rdma_ack_payload_data          (rdma_0_ack_data[42:0]                        ), //i
    .io_rdma_axis_sink_valid           (rdma_0_axis_sink_tvalid                      ), //i
    .io_rdma_axis_sink_ready           (txnEng_io_rdma_axis_sink_ready               ), //o
    .io_rdma_axis_sink_payload_tdata   (rdma_0_axis_sink_tdata[511:0]                ), //i
    .io_rdma_axis_sink_payload_tkeep   (rdma_0_axis_sink_tkeep[63:0]                 ), //i
    .io_rdma_axis_sink_payload_tlast   (rdma_0_axis_sink_tlast                       ), //i
    .io_rdma_axis_src_valid            (txnEng_io_rdma_axis_src_valid                ), //o
    .io_rdma_axis_src_ready            (rdma_0_axis_src_tready                       ), //i
    .io_rdma_axis_src_payload_tdata    (txnEng_io_rdma_axis_src_payload_tdata[511:0] ), //o
    .io_rdma_axis_src_payload_tkeep    (txnEng_io_rdma_axis_src_payload_tkeep[63:0]  ), //o
    .io_rdma_axis_src_payload_tlast    (txnEng_io_rdma_axis_src_payload_tlast        ), //o
    .io_rdmaCtrl_0_en                  (_zz_ctrlR_readRsp_data_6                     ), //i
    .io_rdmaCtrl_0_len                 (_zz_ctrlR_readRsp_data_7[31:0]               ), //i
    .io_rdmaCtrl_0_qpn                 (_zz_ctrlR_readRsp_data_8[9:0]                ), //i
    .io_rdmaCtrl_0_flowId              (_zz_ctrlR_readRsp_data_9[3:0]                ), //i
    .io_rdmaCtrl_1_en                  (_zz_ctrlR_readRsp_data_10                    ), //i
    .io_rdmaCtrl_1_len                 (_zz_ctrlR_readRsp_data_11[31:0]              ), //i
    .io_rdmaCtrl_1_qpn                 (_zz_ctrlR_readRsp_data_12[9:0]               ), //i
    .io_rdmaCtrl_1_flowId              (_zz_ctrlR_readRsp_data_13[3:0]               ), //i
    .io_cntRDMASent                    (txnEng_io_cntRDMASent[31:0]                  ), //o
    .io_cntRDMARecv                    (txnEng_io_cntRDMARecv[31:0]                  ), //o
    .resetn                            (resetn                                       ), //i
    .clk                               (clk                                          )  //i
  );
  assign hostd_bpss_rd_req_valid = hbmHost_io_hostd_bpss_rd_req_valid;
  assign hostd_bpss_rd_req_data = hbmHost_io_hostd_bpss_rd_req_payload_data;
  assign hostd_bpss_wr_req_valid = hbmHost_io_hostd_bpss_wr_req_valid;
  assign hostd_bpss_wr_req_data = hbmHost_io_hostd_bpss_wr_req_payload_data;
  assign hostd_bpss_rd_done_ready = hbmHost_io_hostd_bpss_rd_done_ready;
  assign hostd_bpss_wr_done_ready = hbmHost_io_hostd_bpss_wr_done_ready;
  assign hostd_axis_host_sink_tready = hbmHost_io_hostd_axis_host_sink_ready;
  assign hostd_axis_host_src_tvalid = hbmHost_io_hostd_axis_host_src_valid;
  assign hostd_axis_host_src_tdata = hbmHost_io_hostd_axis_host_src_payload_tdata;
  assign hostd_axis_host_src_tdest = hbmHost_io_hostd_axis_host_src_payload_tdest;
  assign hostd_axis_host_src_tkeep = hbmHost_io_hostd_axis_host_src_payload_tkeep;
  assign hostd_axis_host_src_tlast = hbmHost_io_hostd_axis_host_src_payload_tlast;
  assign axi_mem_0_awvalid = hbmHost_io_axi_cmem_aw_valid;
  assign axi_mem_0_awaddr = hbmHost_io_axi_cmem_aw_payload_addr;
  assign axi_mem_0_awid = hbmHost_io_axi_cmem_aw_payload_id;
  assign axi_mem_0_awlen = hbmHost_io_axi_cmem_aw_payload_len;
  assign axi_mem_0_awsize = hbmHost_io_axi_cmem_aw_payload_size;
  assign axi_mem_0_awburst = hbmHost_io_axi_cmem_aw_payload_burst;
  assign axi_mem_0_wvalid = hbmHost_io_axi_cmem_w_valid;
  assign axi_mem_0_wdata = hbmHost_io_axi_cmem_w_payload_data;
  assign axi_mem_0_wstrb = hbmHost_io_axi_cmem_w_payload_strb;
  assign axi_mem_0_wlast = hbmHost_io_axi_cmem_w_payload_last;
  assign axi_mem_0_bready = hbmHost_io_axi_cmem_b_ready;
  assign axi_mem_0_arvalid = hbmHost_io_axi_cmem_ar_valid;
  assign axi_mem_0_araddr = hbmHost_io_axi_cmem_ar_payload_addr;
  assign axi_mem_0_arid = hbmHost_io_axi_cmem_ar_payload_id;
  assign axi_mem_0_arlen = hbmHost_io_axi_cmem_ar_payload_len;
  assign axi_mem_0_arsize = hbmHost_io_axi_cmem_ar_payload_size;
  assign axi_mem_0_arburst = hbmHost_io_axi_cmem_ar_payload_burst;
  assign axi_mem_0_rready = hbmHost_io_axi_cmem_r_ready;
  assign axi_mem_1_awvalid = txnEng_io_node_axi_0_aw_valid;
  assign axi_mem_1_awaddr = txnEng_io_node_axi_0_aw_payload_addr;
  assign axi_mem_1_awid = txnEng_io_node_axi_0_aw_payload_id;
  assign axi_mem_1_awlen = txnEng_io_node_axi_0_aw_payload_len;
  assign axi_mem_1_awsize = txnEng_io_node_axi_0_aw_payload_size;
  assign axi_mem_1_awburst = txnEng_io_node_axi_0_aw_payload_burst;
  assign axi_mem_1_wvalid = txnEng_io_node_axi_0_w_valid;
  assign axi_mem_1_wdata = txnEng_io_node_axi_0_w_payload_data;
  assign axi_mem_1_wstrb = txnEng_io_node_axi_0_w_payload_strb;
  assign axi_mem_1_wlast = txnEng_io_node_axi_0_w_payload_last;
  assign axi_mem_1_bready = txnEng_io_node_axi_0_b_ready;
  assign axi_mem_1_arvalid = txnEng_io_node_axi_0_ar_valid;
  assign axi_mem_1_araddr = txnEng_io_node_axi_0_ar_payload_addr;
  assign axi_mem_1_arid = txnEng_io_node_axi_0_ar_payload_id;
  assign axi_mem_1_arlen = txnEng_io_node_axi_0_ar_payload_len;
  assign axi_mem_1_arsize = txnEng_io_node_axi_0_ar_payload_size;
  assign axi_mem_1_arburst = txnEng_io_node_axi_0_ar_payload_burst;
  assign axi_mem_1_rready = txnEng_io_node_axi_0_r_ready;
  assign axi_mem_2_awvalid = txnEng_io_node_axi_1_aw_valid;
  assign axi_mem_2_awaddr = txnEng_io_node_axi_1_aw_payload_addr;
  assign axi_mem_2_awid = txnEng_io_node_axi_1_aw_payload_id;
  assign axi_mem_2_awlen = txnEng_io_node_axi_1_aw_payload_len;
  assign axi_mem_2_awsize = txnEng_io_node_axi_1_aw_payload_size;
  assign axi_mem_2_awburst = txnEng_io_node_axi_1_aw_payload_burst;
  assign axi_mem_2_wvalid = txnEng_io_node_axi_1_w_valid;
  assign axi_mem_2_wdata = txnEng_io_node_axi_1_w_payload_data;
  assign axi_mem_2_wstrb = txnEng_io_node_axi_1_w_payload_strb;
  assign axi_mem_2_wlast = txnEng_io_node_axi_1_w_payload_last;
  assign axi_mem_2_bready = txnEng_io_node_axi_1_b_ready;
  assign axi_mem_2_arvalid = txnEng_io_node_axi_1_ar_valid;
  assign axi_mem_2_araddr = txnEng_io_node_axi_1_ar_payload_addr;
  assign axi_mem_2_arid = txnEng_io_node_axi_1_ar_payload_id;
  assign axi_mem_2_arlen = txnEng_io_node_axi_1_ar_payload_len;
  assign axi_mem_2_arsize = txnEng_io_node_axi_1_ar_payload_size;
  assign axi_mem_2_arburst = txnEng_io_node_axi_1_ar_payload_burst;
  assign axi_mem_2_rready = txnEng_io_node_axi_1_r_ready;
  assign axi_mem_3_awvalid = txnEng_io_node_cmdAxi_0_aw_valid;
  assign axi_mem_3_awaddr = txnEng_io_node_cmdAxi_0_aw_payload_addr;
  assign axi_mem_3_awid = txnEng_io_node_cmdAxi_0_aw_payload_id;
  assign axi_mem_3_awlen = txnEng_io_node_cmdAxi_0_aw_payload_len;
  assign axi_mem_3_awsize = txnEng_io_node_cmdAxi_0_aw_payload_size;
  assign axi_mem_3_awburst = txnEng_io_node_cmdAxi_0_aw_payload_burst;
  assign axi_mem_3_wvalid = txnEng_io_node_cmdAxi_0_w_valid;
  assign axi_mem_3_wdata = txnEng_io_node_cmdAxi_0_w_payload_data;
  assign axi_mem_3_wstrb = txnEng_io_node_cmdAxi_0_w_payload_strb;
  assign axi_mem_3_wlast = txnEng_io_node_cmdAxi_0_w_payload_last;
  assign axi_mem_3_bready = txnEng_io_node_cmdAxi_0_b_ready;
  assign axi_mem_3_arvalid = txnEng_io_node_cmdAxi_0_ar_valid;
  assign axi_mem_3_araddr = txnEng_io_node_cmdAxi_0_ar_payload_addr;
  assign axi_mem_3_arid = txnEng_io_node_cmdAxi_0_ar_payload_id;
  assign axi_mem_3_arlen = txnEng_io_node_cmdAxi_0_ar_payload_len;
  assign axi_mem_3_arsize = txnEng_io_node_cmdAxi_0_ar_payload_size;
  assign axi_mem_3_arburst = txnEng_io_node_cmdAxi_0_ar_payload_burst;
  assign axi_mem_3_rready = txnEng_io_node_cmdAxi_0_r_ready;
  assign rdma_0_rd_req_ready = txnEng_io_rdma_rd_req_ready;
  assign rdma_0_wr_req_ready = txnEng_io_rdma_wr_req_ready;
  assign rdma_0_sq_valid = txnEng_io_rdma_sq_valid;
  assign rdma_0_sq_data = txnEng_io_rdma_sq_payload_data;
  assign rdma_0_ack_ready = txnEng_io_rdma_ack_ready;
  assign rdma_0_axis_sink_tready = txnEng_io_rdma_axis_sink_ready;
  assign rdma_0_axis_src_tvalid = txnEng_io_rdma_axis_src_valid;
  assign rdma_0_axis_src_tdata = txnEng_io_rdma_axis_src_payload_tdata;
  assign rdma_0_axis_src_tkeep = txnEng_io_rdma_axis_src_payload_tkeep;
  assign rdma_0_axis_src_tlast = txnEng_io_rdma_axis_src_payload_tlast;
  assign ctrlR_readHaltRequest = 1'b0;
  assign ctrlR_writeHaltRequest = 1'b0;
  assign ctrlR_writeJoinEvent_fire = (ctrlR_writeJoinEvent_valid && ctrlR_writeJoinEvent_ready);
  assign ctrlR_writeJoinEvent_valid = (axi_ctrl_awvalid && axi_ctrl_wvalid);
  assign axi_ctrl_awready = ctrlR_writeJoinEvent_fire;
  assign axi_ctrl_wready = ctrlR_writeJoinEvent_fire;
  assign ctrlR_writeJoinEvent_translated_valid = ctrlR_writeJoinEvent_valid;
  assign ctrlR_writeJoinEvent_ready = ctrlR_writeJoinEvent_translated_ready;
  assign ctrlR_writeJoinEvent_translated_payload_resp = ctrlR_writeRsp_resp;
  assign _zz_axi_ctrl_bvalid = (! ctrlR_writeHaltRequest);
  assign ctrlR_writeJoinEvent_translated_ready = (_zz_ctrlR_writeJoinEvent_translated_ready && _zz_axi_ctrl_bvalid);
  always @(*) begin
    _zz_ctrlR_writeJoinEvent_translated_ready = axi_ctrl_bready;
    if(when_Stream_l368) begin
      _zz_ctrlR_writeJoinEvent_translated_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! _zz_axi_ctrl_bvalid_1);
  assign _zz_axi_ctrl_bvalid_1 = _zz_axi_ctrl_bvalid_2;
  assign axi_ctrl_bvalid = _zz_axi_ctrl_bvalid_1;
  assign axi_ctrl_bresp = _zz_axi_ctrl_bresp;
  always @(*) begin
    axi_ctrl_arready = ctrlR_readDataStage_ready;
    if(when_Stream_l368_1) begin
      axi_ctrl_arready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! ctrlR_readDataStage_valid);
  assign ctrlR_readDataStage_valid = axi_ctrl_ar_rValid;
  assign ctrlR_readDataStage_payload_addr = axi_ctrl_ar_rData_addr;
  assign ctrlR_readDataStage_payload_prot = axi_ctrl_ar_rData_prot;
  assign _zz_axi_ctrl_rvalid = (! ctrlR_readHaltRequest);
  assign ctrlR_readDataStage_ready = (axi_ctrl_rready && _zz_axi_ctrl_rvalid);
  assign axi_ctrl_rvalid = (ctrlR_readDataStage_valid && _zz_axi_ctrl_rvalid);
  assign axi_ctrl_rdata = ctrlR_readRsp_data;
  assign axi_ctrl_rresp = ctrlR_readRsp_resp;
  assign ctrlR_writeRsp_resp = 2'b00;
  assign ctrlR_readRsp_resp = 2'b00;
  always @(*) begin
    ctrlR_readRsp_data = 64'h0;
    case(ctrlR_readAddressMasked)
      64'h0 : begin
        ctrlR_readRsp_data[1 : 0] = _zz_ctrlR_readRsp_data;
      end
      64'h0000000000000008 : begin
        ctrlR_readRsp_data[63 : 0] = _zz_ctrlR_readRsp_data_1;
      end
      64'h0000000000000010 : begin
        ctrlR_readRsp_data[63 : 0] = _zz_ctrlR_readRsp_data_2;
      end
      64'h0000000000000018 : begin
        ctrlR_readRsp_data[15 : 0] = _zz_ctrlR_readRsp_data_3;
      end
      64'h0000000000000020 : begin
        ctrlR_readRsp_data[63 : 0] = _zz_ctrlR_readRsp_data_4;
      end
      64'h0000000000000028 : begin
        ctrlR_readRsp_data[5 : 0] = _zz_ctrlR_readRsp_data_5;
      end
      64'h0000000000000030 : begin
        ctrlR_readRsp_data[63 : 0] = hbmHost_io_cntDone;
      end
      64'h0000000000000038 : begin
        ctrlR_readRsp_data[0 : 0] = _zz_ctrlR_readRsp_data_6;
        ctrlR_readRsp_data[32 : 1] = _zz_ctrlR_readRsp_data_7;
        ctrlR_readRsp_data[42 : 33] = _zz_ctrlR_readRsp_data_8;
        ctrlR_readRsp_data[60 : 57] = _zz_ctrlR_readRsp_data_9;
      end
      64'h0000000000000040 : begin
        ctrlR_readRsp_data[0 : 0] = _zz_ctrlR_readRsp_data_10;
        ctrlR_readRsp_data[32 : 1] = _zz_ctrlR_readRsp_data_11;
        ctrlR_readRsp_data[42 : 33] = _zz_ctrlR_readRsp_data_12;
        ctrlR_readRsp_data[60 : 57] = _zz_ctrlR_readRsp_data_13;
      end
      64'h0000000000000048 : begin
        ctrlR_readRsp_data[0 : 0] = when_Types_l284;
      end
      64'h0000000000000050 : begin
        ctrlR_readRsp_data[0 : 0] = _zz_ctrlR_readRsp_data_14;
      end
      64'h0000000000000058 : begin
        ctrlR_readRsp_data[31 : 0] = _zz_ctrlR_readRsp_data_15;
      end
      64'h0000000000000060 : begin
        ctrlR_readRsp_data[31 : 0] = _zz_ctrlR_readRsp_data_16;
      end
      64'h0000000000000068 : begin
        ctrlR_readRsp_data[0 : 0] = txnEng_io_node_done_0;
      end
      64'h0000000000000070 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntClk_0;
      end
      64'h0000000000000078 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntTxnLd_0;
      end
      64'h0000000000000080 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntTxnCmt_0;
      end
      64'h0000000000000088 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntTxnAbt_0;
      end
      64'h0000000000000090 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntLockLoc_0;
      end
      64'h0000000000000098 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntLockRmt_0;
      end
      64'h00000000000000a0 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntLockDenyLoc_0;
      end
      64'h00000000000000a8 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_node_cntLockDenyRmt_0;
      end
      64'h00000000000000b0 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_cntRDMASent;
      end
      64'h00000000000000b8 : begin
        ctrlR_readRsp_data[31 : 0] = txnEng_io_cntRDMARecv;
      end
      default : begin
      end
    endcase
  end

  assign ctrlR_readAddressMasked = (ctrlR_readDataStage_payload_addr & (~ 64'h0000000000000007));
  assign ctrlR_writeAddressMasked = (axi_ctrl_awaddr & (~ 64'h0000000000000007));
  assign ctrlR_writeOccur = (ctrlR_writeJoinEvent_valid && ctrlR_writeJoinEvent_ready);
  assign ctrlR_readOccur = (axi_ctrl_rvalid && axi_ctrl_rready);
  assign when_Types_l264 = (|_zz_ctrlR_readRsp_data);
  assign when_BusSlaveFactory_l962 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_1 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_2 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_3 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_4 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_5 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_6 = axi_ctrl_wstrb[5];
  assign when_BusSlaveFactory_l962_7 = axi_ctrl_wstrb[6];
  assign when_BusSlaveFactory_l962_8 = axi_ctrl_wstrb[7];
  assign when_BusSlaveFactory_l962_9 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_10 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_11 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_12 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_13 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_14 = axi_ctrl_wstrb[5];
  assign when_BusSlaveFactory_l962_15 = axi_ctrl_wstrb[6];
  assign when_BusSlaveFactory_l962_16 = axi_ctrl_wstrb[7];
  assign when_BusSlaveFactory_l962_17 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_18 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_19 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_20 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_21 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_22 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_23 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_24 = axi_ctrl_wstrb[5];
  assign when_BusSlaveFactory_l962_25 = axi_ctrl_wstrb[6];
  assign when_BusSlaveFactory_l962_26 = axi_ctrl_wstrb[7];
  assign when_BusSlaveFactory_l962_27 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_28 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_29 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_30 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_31 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_32 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_33 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_34 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_35 = axi_ctrl_wstrb[5];
  assign when_BusSlaveFactory_l962_36 = axi_ctrl_wstrb[7];
  assign when_BusSlaveFactory_l962_37 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_38 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_39 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_40 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_41 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_42 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_43 = axi_ctrl_wstrb[4];
  assign when_BusSlaveFactory_l962_44 = axi_ctrl_wstrb[5];
  assign when_BusSlaveFactory_l962_45 = axi_ctrl_wstrb[7];
  assign when_BusSlaveFactory_l962_46 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_47 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_48 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_49 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_50 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_51 = axi_ctrl_wstrb[3];
  assign when_BusSlaveFactory_l962_52 = axi_ctrl_wstrb[0];
  assign when_BusSlaveFactory_l962_53 = axi_ctrl_wstrb[1];
  assign when_BusSlaveFactory_l962_54 = axi_ctrl_wstrb[2];
  assign when_BusSlaveFactory_l962_55 = axi_ctrl_wstrb[3];
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_axi_ctrl_bvalid_2 <= 1'b0;
      axi_ctrl_ar_rValid <= 1'b0;
    end else begin
      if(_zz_ctrlR_writeJoinEvent_translated_ready) begin
        _zz_axi_ctrl_bvalid_2 <= (ctrlR_writeJoinEvent_translated_valid && _zz_axi_ctrl_bvalid);
      end
      if(axi_ctrl_arready) begin
        axi_ctrl_ar_rValid <= axi_ctrl_arvalid;
      end
    end
  end

  always @(posedge clk) begin
    if(_zz_ctrlR_writeJoinEvent_translated_ready) begin
      _zz_axi_ctrl_bresp <= ctrlR_writeJoinEvent_translated_payload_resp;
    end
    if(axi_ctrl_arready) begin
      axi_ctrl_ar_rData_addr <= axi_ctrl_araddr;
      axi_ctrl_ar_rData_prot <= axi_ctrl_arprot;
    end
    if(when_Types_l264) begin
      _zz_ctrlR_readRsp_data <= 2'b00;
    end
    if(when_Types_l284) begin
      when_Types_l284 <= 1'b0;
    end
    case(ctrlR_writeAddressMasked)
      64'h0 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962) begin
            _zz_ctrlR_readRsp_data[1 : 0] <= axi_ctrl_wdata[1 : 0];
          end
        end
      end
      64'h0000000000000008 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_1) begin
            _zz_ctrlR_readRsp_data_1[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_2) begin
            _zz_ctrlR_readRsp_data_1[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_3) begin
            _zz_ctrlR_readRsp_data_1[23 : 16] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_4) begin
            _zz_ctrlR_readRsp_data_1[31 : 24] <= axi_ctrl_wdata[31 : 24];
          end
          if(when_BusSlaveFactory_l962_5) begin
            _zz_ctrlR_readRsp_data_1[39 : 32] <= axi_ctrl_wdata[39 : 32];
          end
          if(when_BusSlaveFactory_l962_6) begin
            _zz_ctrlR_readRsp_data_1[47 : 40] <= axi_ctrl_wdata[47 : 40];
          end
          if(when_BusSlaveFactory_l962_7) begin
            _zz_ctrlR_readRsp_data_1[55 : 48] <= axi_ctrl_wdata[55 : 48];
          end
          if(when_BusSlaveFactory_l962_8) begin
            _zz_ctrlR_readRsp_data_1[63 : 56] <= axi_ctrl_wdata[63 : 56];
          end
        end
      end
      64'h0000000000000010 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_9) begin
            _zz_ctrlR_readRsp_data_2[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_10) begin
            _zz_ctrlR_readRsp_data_2[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_11) begin
            _zz_ctrlR_readRsp_data_2[23 : 16] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_12) begin
            _zz_ctrlR_readRsp_data_2[31 : 24] <= axi_ctrl_wdata[31 : 24];
          end
          if(when_BusSlaveFactory_l962_13) begin
            _zz_ctrlR_readRsp_data_2[39 : 32] <= axi_ctrl_wdata[39 : 32];
          end
          if(when_BusSlaveFactory_l962_14) begin
            _zz_ctrlR_readRsp_data_2[47 : 40] <= axi_ctrl_wdata[47 : 40];
          end
          if(when_BusSlaveFactory_l962_15) begin
            _zz_ctrlR_readRsp_data_2[55 : 48] <= axi_ctrl_wdata[55 : 48];
          end
          if(when_BusSlaveFactory_l962_16) begin
            _zz_ctrlR_readRsp_data_2[63 : 56] <= axi_ctrl_wdata[63 : 56];
          end
        end
      end
      64'h0000000000000018 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_17) begin
            _zz_ctrlR_readRsp_data_3[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_18) begin
            _zz_ctrlR_readRsp_data_3[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
        end
      end
      64'h0000000000000020 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_19) begin
            _zz_ctrlR_readRsp_data_4[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_20) begin
            _zz_ctrlR_readRsp_data_4[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_21) begin
            _zz_ctrlR_readRsp_data_4[23 : 16] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_22) begin
            _zz_ctrlR_readRsp_data_4[31 : 24] <= axi_ctrl_wdata[31 : 24];
          end
          if(when_BusSlaveFactory_l962_23) begin
            _zz_ctrlR_readRsp_data_4[39 : 32] <= axi_ctrl_wdata[39 : 32];
          end
          if(when_BusSlaveFactory_l962_24) begin
            _zz_ctrlR_readRsp_data_4[47 : 40] <= axi_ctrl_wdata[47 : 40];
          end
          if(when_BusSlaveFactory_l962_25) begin
            _zz_ctrlR_readRsp_data_4[55 : 48] <= axi_ctrl_wdata[55 : 48];
          end
          if(when_BusSlaveFactory_l962_26) begin
            _zz_ctrlR_readRsp_data_4[63 : 56] <= axi_ctrl_wdata[63 : 56];
          end
        end
      end
      64'h0000000000000028 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_27) begin
            _zz_ctrlR_readRsp_data_5[5 : 0] <= axi_ctrl_wdata[5 : 0];
          end
        end
      end
      64'h0000000000000038 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_28) begin
            _zz_ctrlR_readRsp_data_6 <= axi_ctrl_wdata[0];
          end
          if(when_BusSlaveFactory_l962_29) begin
            _zz_ctrlR_readRsp_data_7[6 : 0] <= axi_ctrl_wdata[7 : 1];
          end
          if(when_BusSlaveFactory_l962_30) begin
            _zz_ctrlR_readRsp_data_7[14 : 7] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_31) begin
            _zz_ctrlR_readRsp_data_7[22 : 15] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_32) begin
            _zz_ctrlR_readRsp_data_7[30 : 23] <= axi_ctrl_wdata[31 : 24];
          end
          if(when_BusSlaveFactory_l962_33) begin
            _zz_ctrlR_readRsp_data_7[31 : 31] <= axi_ctrl_wdata[32 : 32];
          end
          if(when_BusSlaveFactory_l962_34) begin
            _zz_ctrlR_readRsp_data_8[6 : 0] <= axi_ctrl_wdata[39 : 33];
          end
          if(when_BusSlaveFactory_l962_35) begin
            _zz_ctrlR_readRsp_data_8[9 : 7] <= axi_ctrl_wdata[42 : 40];
          end
          if(when_BusSlaveFactory_l962_36) begin
            _zz_ctrlR_readRsp_data_9[3 : 0] <= axi_ctrl_wdata[60 : 57];
          end
        end
      end
      64'h0000000000000040 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_37) begin
            _zz_ctrlR_readRsp_data_10 <= axi_ctrl_wdata[0];
          end
          if(when_BusSlaveFactory_l962_38) begin
            _zz_ctrlR_readRsp_data_11[6 : 0] <= axi_ctrl_wdata[7 : 1];
          end
          if(when_BusSlaveFactory_l962_39) begin
            _zz_ctrlR_readRsp_data_11[14 : 7] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_40) begin
            _zz_ctrlR_readRsp_data_11[22 : 15] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_41) begin
            _zz_ctrlR_readRsp_data_11[30 : 23] <= axi_ctrl_wdata[31 : 24];
          end
          if(when_BusSlaveFactory_l962_42) begin
            _zz_ctrlR_readRsp_data_11[31 : 31] <= axi_ctrl_wdata[32 : 32];
          end
          if(when_BusSlaveFactory_l962_43) begin
            _zz_ctrlR_readRsp_data_12[6 : 0] <= axi_ctrl_wdata[39 : 33];
          end
          if(when_BusSlaveFactory_l962_44) begin
            _zz_ctrlR_readRsp_data_12[9 : 7] <= axi_ctrl_wdata[42 : 40];
          end
          if(when_BusSlaveFactory_l962_45) begin
            _zz_ctrlR_readRsp_data_13[3 : 0] <= axi_ctrl_wdata[60 : 57];
          end
        end
      end
      64'h0000000000000048 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_46) begin
            when_Types_l284 <= axi_ctrl_wdata[0];
          end
        end
      end
      64'h0000000000000050 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_47) begin
            _zz_ctrlR_readRsp_data_14[0 : 0] <= axi_ctrl_wdata[0 : 0];
          end
        end
      end
      64'h0000000000000058 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_48) begin
            _zz_ctrlR_readRsp_data_15[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_49) begin
            _zz_ctrlR_readRsp_data_15[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_50) begin
            _zz_ctrlR_readRsp_data_15[23 : 16] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_51) begin
            _zz_ctrlR_readRsp_data_15[31 : 24] <= axi_ctrl_wdata[31 : 24];
          end
        end
      end
      64'h0000000000000060 : begin
        if(ctrlR_writeOccur) begin
          if(when_BusSlaveFactory_l962_52) begin
            _zz_ctrlR_readRsp_data_16[7 : 0] <= axi_ctrl_wdata[7 : 0];
          end
          if(when_BusSlaveFactory_l962_53) begin
            _zz_ctrlR_readRsp_data_16[15 : 8] <= axi_ctrl_wdata[15 : 8];
          end
          if(when_BusSlaveFactory_l962_54) begin
            _zz_ctrlR_readRsp_data_16[23 : 16] <= axi_ctrl_wdata[23 : 16];
          end
          if(when_BusSlaveFactory_l962_55) begin
            _zz_ctrlR_readRsp_data_16[31 : 24] <= axi_ctrl_wdata[31 : 24];
          end
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module WrapNodeNet (
  output              io_node_axi_0_aw_valid,
  input               io_node_axi_0_aw_ready,
  output     [63:0]   io_node_axi_0_aw_payload_addr,
  output     [5:0]    io_node_axi_0_aw_payload_id,
  output     [7:0]    io_node_axi_0_aw_payload_len,
  output     [2:0]    io_node_axi_0_aw_payload_size,
  output     [1:0]    io_node_axi_0_aw_payload_burst,
  output              io_node_axi_0_w_valid,
  input               io_node_axi_0_w_ready,
  output     [511:0]  io_node_axi_0_w_payload_data,
  output     [63:0]   io_node_axi_0_w_payload_strb,
  output              io_node_axi_0_w_payload_last,
  input               io_node_axi_0_b_valid,
  output              io_node_axi_0_b_ready,
  input      [5:0]    io_node_axi_0_b_payload_id,
  input      [1:0]    io_node_axi_0_b_payload_resp,
  output              io_node_axi_0_ar_valid,
  input               io_node_axi_0_ar_ready,
  output     [63:0]   io_node_axi_0_ar_payload_addr,
  output     [5:0]    io_node_axi_0_ar_payload_id,
  output     [7:0]    io_node_axi_0_ar_payload_len,
  output     [2:0]    io_node_axi_0_ar_payload_size,
  output     [1:0]    io_node_axi_0_ar_payload_burst,
  input               io_node_axi_0_r_valid,
  output              io_node_axi_0_r_ready,
  input      [511:0]  io_node_axi_0_r_payload_data,
  input      [5:0]    io_node_axi_0_r_payload_id,
  input      [1:0]    io_node_axi_0_r_payload_resp,
  input               io_node_axi_0_r_payload_last,
  output              io_node_axi_1_aw_valid,
  input               io_node_axi_1_aw_ready,
  output     [63:0]   io_node_axi_1_aw_payload_addr,
  output     [5:0]    io_node_axi_1_aw_payload_id,
  output     [7:0]    io_node_axi_1_aw_payload_len,
  output     [2:0]    io_node_axi_1_aw_payload_size,
  output     [1:0]    io_node_axi_1_aw_payload_burst,
  output              io_node_axi_1_w_valid,
  input               io_node_axi_1_w_ready,
  output     [511:0]  io_node_axi_1_w_payload_data,
  output     [63:0]   io_node_axi_1_w_payload_strb,
  output              io_node_axi_1_w_payload_last,
  input               io_node_axi_1_b_valid,
  output              io_node_axi_1_b_ready,
  input      [5:0]    io_node_axi_1_b_payload_id,
  input      [1:0]    io_node_axi_1_b_payload_resp,
  output              io_node_axi_1_ar_valid,
  input               io_node_axi_1_ar_ready,
  output     [63:0]   io_node_axi_1_ar_payload_addr,
  output     [5:0]    io_node_axi_1_ar_payload_id,
  output     [7:0]    io_node_axi_1_ar_payload_len,
  output     [2:0]    io_node_axi_1_ar_payload_size,
  output     [1:0]    io_node_axi_1_ar_payload_burst,
  input               io_node_axi_1_r_valid,
  output              io_node_axi_1_r_ready,
  input      [511:0]  io_node_axi_1_r_payload_data,
  input      [5:0]    io_node_axi_1_r_payload_id,
  input      [1:0]    io_node_axi_1_r_payload_resp,
  input               io_node_axi_1_r_payload_last,
  output              io_node_cmdAxi_0_aw_valid,
  input               io_node_cmdAxi_0_aw_ready,
  output     [63:0]   io_node_cmdAxi_0_aw_payload_addr,
  output     [5:0]    io_node_cmdAxi_0_aw_payload_id,
  output     [7:0]    io_node_cmdAxi_0_aw_payload_len,
  output     [2:0]    io_node_cmdAxi_0_aw_payload_size,
  output     [1:0]    io_node_cmdAxi_0_aw_payload_burst,
  output              io_node_cmdAxi_0_w_valid,
  input               io_node_cmdAxi_0_w_ready,
  output     [511:0]  io_node_cmdAxi_0_w_payload_data,
  output     [63:0]   io_node_cmdAxi_0_w_payload_strb,
  output              io_node_cmdAxi_0_w_payload_last,
  input               io_node_cmdAxi_0_b_valid,
  output              io_node_cmdAxi_0_b_ready,
  input      [5:0]    io_node_cmdAxi_0_b_payload_id,
  input      [1:0]    io_node_cmdAxi_0_b_payload_resp,
  output              io_node_cmdAxi_0_ar_valid,
  input               io_node_cmdAxi_0_ar_ready,
  output     [63:0]   io_node_cmdAxi_0_ar_payload_addr,
  output     [5:0]    io_node_cmdAxi_0_ar_payload_id,
  output     [7:0]    io_node_cmdAxi_0_ar_payload_len,
  output     [2:0]    io_node_cmdAxi_0_ar_payload_size,
  output     [1:0]    io_node_cmdAxi_0_ar_payload_burst,
  input               io_node_cmdAxi_0_r_valid,
  output              io_node_cmdAxi_0_r_ready,
  input      [511:0]  io_node_cmdAxi_0_r_payload_data,
  input      [5:0]    io_node_cmdAxi_0_r_payload_id,
  input      [1:0]    io_node_cmdAxi_0_r_payload_resp,
  input               io_node_cmdAxi_0_r_payload_last,
  input      [0:0]    io_node_nodeId,
  input      [31:0]   io_node_txnNumTotal,
  input      [31:0]   io_node_cmdAddrOffs_0,
  input               io_node_start,
  output              io_node_done_0,
  output     [31:0]   io_node_cntTxnCmt_0,
  output     [31:0]   io_node_cntTxnAbt_0,
  output     [31:0]   io_node_cntTxnLd_0,
  output     [31:0]   io_node_cntLockLoc_0,
  output     [31:0]   io_node_cntLockRmt_0,
  output     [31:0]   io_node_cntLockDenyLoc_0,
  output     [31:0]   io_node_cntLockDenyRmt_0,
  output     [31:0]   io_node_cntClk_0,
  input               io_rdma_rd_req_valid,
  output              io_rdma_rd_req_ready,
  input      [95:0]   io_rdma_rd_req_payload_data,
  input               io_rdma_wr_req_valid,
  output              io_rdma_wr_req_ready,
  input      [95:0]   io_rdma_wr_req_payload_data,
  output              io_rdma_sq_valid,
  input               io_rdma_sq_ready,
  output     [543:0]  io_rdma_sq_payload_data,
  input               io_rdma_ack_valid,
  output              io_rdma_ack_ready,
  input      [42:0]   io_rdma_ack_payload_data,
  input               io_rdma_axis_sink_valid,
  output              io_rdma_axis_sink_ready,
  input      [511:0]  io_rdma_axis_sink_payload_tdata,
  input      [63:0]   io_rdma_axis_sink_payload_tkeep,
  input               io_rdma_axis_sink_payload_tlast,
  output              io_rdma_axis_src_valid,
  input               io_rdma_axis_src_ready,
  output     [511:0]  io_rdma_axis_src_payload_tdata,
  output     [63:0]   io_rdma_axis_src_payload_tkeep,
  output              io_rdma_axis_src_payload_tlast,
  input               io_rdmaCtrl_0_en,
  input      [31:0]   io_rdmaCtrl_0_len,
  input      [9:0]    io_rdmaCtrl_0_qpn,
  input      [3:0]    io_rdmaCtrl_0_flowId,
  input               io_rdmaCtrl_1_en,
  input      [31:0]   io_rdmaCtrl_1_len,
  input      [9:0]    io_rdmaCtrl_1_qpn,
  input      [3:0]    io_rdmaCtrl_1_flowId,
  output     [31:0]   io_cntRDMASent,
  output     [31:0]   io_cntRDMARecv,
  input               resetn,
  input               clk
);

  wire                nodeFlow_io_axi_0_ar_valid;
  wire       [63:0]   nodeFlow_io_axi_0_ar_payload_addr;
  wire       [5:0]    nodeFlow_io_axi_0_ar_payload_id;
  wire       [7:0]    nodeFlow_io_axi_0_ar_payload_len;
  wire       [2:0]    nodeFlow_io_axi_0_ar_payload_size;
  wire       [1:0]    nodeFlow_io_axi_0_ar_payload_burst;
  wire                nodeFlow_io_axi_0_aw_valid;
  wire       [63:0]   nodeFlow_io_axi_0_aw_payload_addr;
  wire       [5:0]    nodeFlow_io_axi_0_aw_payload_id;
  wire       [7:0]    nodeFlow_io_axi_0_aw_payload_len;
  wire       [2:0]    nodeFlow_io_axi_0_aw_payload_size;
  wire       [1:0]    nodeFlow_io_axi_0_aw_payload_burst;
  wire                nodeFlow_io_axi_0_w_valid;
  wire       [511:0]  nodeFlow_io_axi_0_w_payload_data;
  wire       [63:0]   nodeFlow_io_axi_0_w_payload_strb;
  wire                nodeFlow_io_axi_0_w_payload_last;
  wire                nodeFlow_io_axi_0_r_ready;
  wire                nodeFlow_io_axi_0_b_ready;
  wire                nodeFlow_io_axi_1_ar_valid;
  wire       [63:0]   nodeFlow_io_axi_1_ar_payload_addr;
  wire       [5:0]    nodeFlow_io_axi_1_ar_payload_id;
  wire       [7:0]    nodeFlow_io_axi_1_ar_payload_len;
  wire       [2:0]    nodeFlow_io_axi_1_ar_payload_size;
  wire       [1:0]    nodeFlow_io_axi_1_ar_payload_burst;
  wire                nodeFlow_io_axi_1_aw_valid;
  wire       [63:0]   nodeFlow_io_axi_1_aw_payload_addr;
  wire       [5:0]    nodeFlow_io_axi_1_aw_payload_id;
  wire       [7:0]    nodeFlow_io_axi_1_aw_payload_len;
  wire       [2:0]    nodeFlow_io_axi_1_aw_payload_size;
  wire       [1:0]    nodeFlow_io_axi_1_aw_payload_burst;
  wire                nodeFlow_io_axi_1_w_valid;
  wire       [511:0]  nodeFlow_io_axi_1_w_payload_data;
  wire       [63:0]   nodeFlow_io_axi_1_w_payload_strb;
  wire                nodeFlow_io_axi_1_w_payload_last;
  wire                nodeFlow_io_axi_1_r_ready;
  wire                nodeFlow_io_axi_1_b_ready;
  wire                nodeFlow_io_cmdAxi_0_ar_valid;
  wire       [63:0]   nodeFlow_io_cmdAxi_0_ar_payload_addr;
  wire       [5:0]    nodeFlow_io_cmdAxi_0_ar_payload_id;
  wire       [7:0]    nodeFlow_io_cmdAxi_0_ar_payload_len;
  wire       [2:0]    nodeFlow_io_cmdAxi_0_ar_payload_size;
  wire       [1:0]    nodeFlow_io_cmdAxi_0_ar_payload_burst;
  wire                nodeFlow_io_cmdAxi_0_aw_valid;
  wire       [63:0]   nodeFlow_io_cmdAxi_0_aw_payload_addr;
  wire       [5:0]    nodeFlow_io_cmdAxi_0_aw_payload_id;
  wire       [7:0]    nodeFlow_io_cmdAxi_0_aw_payload_len;
  wire       [2:0]    nodeFlow_io_cmdAxi_0_aw_payload_size;
  wire       [1:0]    nodeFlow_io_cmdAxi_0_aw_payload_burst;
  wire                nodeFlow_io_cmdAxi_0_w_valid;
  wire       [511:0]  nodeFlow_io_cmdAxi_0_w_payload_data;
  wire       [63:0]   nodeFlow_io_cmdAxi_0_w_payload_strb;
  wire                nodeFlow_io_cmdAxi_0_w_payload_last;
  wire                nodeFlow_io_cmdAxi_0_r_ready;
  wire                nodeFlow_io_cmdAxi_0_b_ready;
  wire                nodeFlow_io_done_0;
  wire       [31:0]   nodeFlow_io_cntTxnCmt_0;
  wire       [31:0]   nodeFlow_io_cntTxnAbt_0;
  wire       [31:0]   nodeFlow_io_cntTxnLd_0;
  wire       [31:0]   nodeFlow_io_cntLockLoc_0;
  wire       [31:0]   nodeFlow_io_cntLockRmt_0;
  wire       [31:0]   nodeFlow_io_cntLockDenyLoc_0;
  wire       [31:0]   nodeFlow_io_cntLockDenyRmt_0;
  wire       [31:0]   nodeFlow_io_cntClk_0;
  wire                nodeFlow_io_sendQ_valid;
  wire       [511:0]  nodeFlow_io_sendQ_payload;
  wire                nodeFlow_io_respQ_valid;
  wire       [511:0]  nodeFlow_io_respQ_payload;
  wire                nodeFlow_io_reqQ_ready;
  wire                nodeFlow_io_recvQ_ready;
  wire                nodeFlow_io_sendStatusVld;
  wire                nodeFlow_io_recvStatusVld;
  wire       [3:0]    nodeFlow_io_nReq;
  wire       [3:0]    nodeFlow_io_nWrCmtReq;
  wire       [3:0]    nodeFlow_io_nRdGetReq;
  wire       [3:0]    nodeFlow_io_nResp;
  wire       [3:0]    nodeFlow_io_nWrCmtResp;
  wire       [3:0]    nodeFlow_io_nRdGetResp;
  wire                rdmaFlowMstr_io_rdma_rd_req_ready;
  wire                rdmaFlowMstr_io_rdma_wr_req_ready;
  wire                rdmaFlowMstr_io_rdma_sq_valid;
  wire       [543:0]  rdmaFlowMstr_io_rdma_sq_payload_data;
  wire                rdmaFlowMstr_io_rdma_ack_ready;
  wire                rdmaFlowMstr_io_rdma_axis_sink_ready;
  wire                rdmaFlowMstr_io_rdma_axis_src_valid;
  wire       [511:0]  rdmaFlowMstr_io_rdma_axis_src_payload_tdata;
  wire       [63:0]   rdmaFlowMstr_io_rdma_axis_src_payload_tkeep;
  wire                rdmaFlowMstr_io_rdma_axis_src_payload_tlast;
  wire                rdmaFlowMstr_io_q_sink_ready;
  wire                rdmaFlowMstr_io_q_src_valid;
  wire       [511:0]  rdmaFlowMstr_io_q_src_payload;
  wire                rdmaFlowSlve_io_rdma_rd_req_ready;
  wire                rdmaFlowSlve_io_rdma_wr_req_ready;
  wire                rdmaFlowSlve_io_rdma_sq_valid;
  wire       [543:0]  rdmaFlowSlve_io_rdma_sq_payload_data;
  wire                rdmaFlowSlve_io_rdma_ack_ready;
  wire                rdmaFlowSlve_io_rdma_axis_sink_ready;
  wire                rdmaFlowSlve_io_rdma_axis_src_valid;
  wire       [511:0]  rdmaFlowSlve_io_rdma_axis_src_payload_tdata;
  wire       [63:0]   rdmaFlowSlve_io_rdma_axis_src_payload_tkeep;
  wire                rdmaFlowSlve_io_rdma_axis_src_payload_tlast;
  wire                rdmaFlowSlve_io_q_sink_ready;
  wire                rdmaFlowSlve_io_q_src_valid;
  wire       [511:0]  rdmaFlowSlve_io_q_src_payload;
  wire                rdmaArb_1_io_rdmaV_0_rd_req_valid;
  wire       [95:0]   rdmaArb_1_io_rdmaV_0_rd_req_payload_data;
  wire                rdmaArb_1_io_rdmaV_0_wr_req_valid;
  wire       [95:0]   rdmaArb_1_io_rdmaV_0_wr_req_payload_data;
  wire                rdmaArb_1_io_rdmaV_0_sq_ready;
  wire                rdmaArb_1_io_rdmaV_0_ack_valid;
  wire       [42:0]   rdmaArb_1_io_rdmaV_0_ack_payload_data;
  wire                rdmaArb_1_io_rdmaV_0_axis_sink_valid;
  wire       [511:0]  rdmaArb_1_io_rdmaV_0_axis_sink_payload_tdata;
  wire       [63:0]   rdmaArb_1_io_rdmaV_0_axis_sink_payload_tkeep;
  wire                rdmaArb_1_io_rdmaV_0_axis_sink_payload_tlast;
  wire                rdmaArb_1_io_rdmaV_0_axis_src_ready;
  wire                rdmaArb_1_io_rdmaV_1_rd_req_valid;
  wire       [95:0]   rdmaArb_1_io_rdmaV_1_rd_req_payload_data;
  wire                rdmaArb_1_io_rdmaV_1_wr_req_valid;
  wire       [95:0]   rdmaArb_1_io_rdmaV_1_wr_req_payload_data;
  wire                rdmaArb_1_io_rdmaV_1_sq_ready;
  wire                rdmaArb_1_io_rdmaV_1_ack_valid;
  wire       [42:0]   rdmaArb_1_io_rdmaV_1_ack_payload_data;
  wire                rdmaArb_1_io_rdmaV_1_axis_sink_valid;
  wire       [511:0]  rdmaArb_1_io_rdmaV_1_axis_sink_payload_tdata;
  wire       [63:0]   rdmaArb_1_io_rdmaV_1_axis_sink_payload_tkeep;
  wire                rdmaArb_1_io_rdmaV_1_axis_sink_payload_tlast;
  wire                rdmaArb_1_io_rdmaV_1_axis_src_ready;
  wire                rdmaArb_1_io_rdmaio_rd_req_ready;
  wire                rdmaArb_1_io_rdmaio_wr_req_ready;
  wire                rdmaArb_1_io_rdmaio_sq_valid;
  wire       [543:0]  rdmaArb_1_io_rdmaio_sq_payload_data;
  wire                rdmaArb_1_io_rdmaio_ack_ready;
  wire                rdmaArb_1_io_rdmaio_axis_sink_ready;
  wire                rdmaArb_1_io_rdmaio_axis_src_valid;
  wire       [511:0]  rdmaArb_1_io_rdmaio_axis_src_payload_tdata;
  wire       [63:0]   rdmaArb_1_io_rdmaio_axis_src_payload_tkeep;
  wire                rdmaArb_1_io_rdmaio_axis_src_payload_tlast;
  wire       [31:0]   _zz_cntSent_valueNext;
  wire       [0:0]    _zz_cntSent_valueNext_1;
  wire       [31:0]   _zz_cntRecv_valueNext;
  wire       [0:0]    _zz_cntRecv_valueNext_1;
  reg                 cntSent_willIncrement;
  reg                 cntSent_willClear;
  reg        [31:0]   cntSent_valueNext;
  reg        [31:0]   cntSent_value;
  wire                cntSent_willOverflowIfInc;
  wire                cntSent_willOverflow;
  reg                 cntRecv_willIncrement;
  reg                 cntRecv_willClear;
  reg        [31:0]   cntRecv_valueNext;
  reg        [31:0]   cntRecv_value;
  wire                cntRecv_willOverflowIfInc;
  wire                cntRecv_willOverflow;
  wire                io_rdma_axis_src_fire;
  wire                io_rdma_axis_sink_fire;
  wire                when_WrapNodeNet_l49;
  wire                when_WrapNodeNet_l52;

  assign _zz_cntSent_valueNext_1 = cntSent_willIncrement;
  assign _zz_cntSent_valueNext = {31'd0, _zz_cntSent_valueNext_1};
  assign _zz_cntRecv_valueNext_1 = cntRecv_willIncrement;
  assign _zz_cntRecv_valueNext = {31'd0, _zz_cntRecv_valueNext_1};
  WrapNode nodeFlow (
    .io_axi_0_aw_valid            (nodeFlow_io_axi_0_aw_valid                ), //o
    .io_axi_0_aw_ready            (io_node_axi_0_aw_ready                    ), //i
    .io_axi_0_aw_payload_addr     (nodeFlow_io_axi_0_aw_payload_addr[63:0]   ), //o
    .io_axi_0_aw_payload_id       (nodeFlow_io_axi_0_aw_payload_id[5:0]      ), //o
    .io_axi_0_aw_payload_len      (nodeFlow_io_axi_0_aw_payload_len[7:0]     ), //o
    .io_axi_0_aw_payload_size     (nodeFlow_io_axi_0_aw_payload_size[2:0]    ), //o
    .io_axi_0_aw_payload_burst    (nodeFlow_io_axi_0_aw_payload_burst[1:0]   ), //o
    .io_axi_0_w_valid             (nodeFlow_io_axi_0_w_valid                 ), //o
    .io_axi_0_w_ready             (io_node_axi_0_w_ready                     ), //i
    .io_axi_0_w_payload_data      (nodeFlow_io_axi_0_w_payload_data[511:0]   ), //o
    .io_axi_0_w_payload_strb      (nodeFlow_io_axi_0_w_payload_strb[63:0]    ), //o
    .io_axi_0_w_payload_last      (nodeFlow_io_axi_0_w_payload_last          ), //o
    .io_axi_0_b_valid             (io_node_axi_0_b_valid                     ), //i
    .io_axi_0_b_ready             (nodeFlow_io_axi_0_b_ready                 ), //o
    .io_axi_0_b_payload_id        (io_node_axi_0_b_payload_id[5:0]           ), //i
    .io_axi_0_b_payload_resp      (io_node_axi_0_b_payload_resp[1:0]         ), //i
    .io_axi_0_ar_valid            (nodeFlow_io_axi_0_ar_valid                ), //o
    .io_axi_0_ar_ready            (io_node_axi_0_ar_ready                    ), //i
    .io_axi_0_ar_payload_addr     (nodeFlow_io_axi_0_ar_payload_addr[63:0]   ), //o
    .io_axi_0_ar_payload_id       (nodeFlow_io_axi_0_ar_payload_id[5:0]      ), //o
    .io_axi_0_ar_payload_len      (nodeFlow_io_axi_0_ar_payload_len[7:0]     ), //o
    .io_axi_0_ar_payload_size     (nodeFlow_io_axi_0_ar_payload_size[2:0]    ), //o
    .io_axi_0_ar_payload_burst    (nodeFlow_io_axi_0_ar_payload_burst[1:0]   ), //o
    .io_axi_0_r_valid             (io_node_axi_0_r_valid                     ), //i
    .io_axi_0_r_ready             (nodeFlow_io_axi_0_r_ready                 ), //o
    .io_axi_0_r_payload_data      (io_node_axi_0_r_payload_data[511:0]       ), //i
    .io_axi_0_r_payload_id        (io_node_axi_0_r_payload_id[5:0]           ), //i
    .io_axi_0_r_payload_resp      (io_node_axi_0_r_payload_resp[1:0]         ), //i
    .io_axi_0_r_payload_last      (io_node_axi_0_r_payload_last              ), //i
    .io_axi_1_aw_valid            (nodeFlow_io_axi_1_aw_valid                ), //o
    .io_axi_1_aw_ready            (io_node_axi_1_aw_ready                    ), //i
    .io_axi_1_aw_payload_addr     (nodeFlow_io_axi_1_aw_payload_addr[63:0]   ), //o
    .io_axi_1_aw_payload_id       (nodeFlow_io_axi_1_aw_payload_id[5:0]      ), //o
    .io_axi_1_aw_payload_len      (nodeFlow_io_axi_1_aw_payload_len[7:0]     ), //o
    .io_axi_1_aw_payload_size     (nodeFlow_io_axi_1_aw_payload_size[2:0]    ), //o
    .io_axi_1_aw_payload_burst    (nodeFlow_io_axi_1_aw_payload_burst[1:0]   ), //o
    .io_axi_1_w_valid             (nodeFlow_io_axi_1_w_valid                 ), //o
    .io_axi_1_w_ready             (io_node_axi_1_w_ready                     ), //i
    .io_axi_1_w_payload_data      (nodeFlow_io_axi_1_w_payload_data[511:0]   ), //o
    .io_axi_1_w_payload_strb      (nodeFlow_io_axi_1_w_payload_strb[63:0]    ), //o
    .io_axi_1_w_payload_last      (nodeFlow_io_axi_1_w_payload_last          ), //o
    .io_axi_1_b_valid             (io_node_axi_1_b_valid                     ), //i
    .io_axi_1_b_ready             (nodeFlow_io_axi_1_b_ready                 ), //o
    .io_axi_1_b_payload_id        (io_node_axi_1_b_payload_id[5:0]           ), //i
    .io_axi_1_b_payload_resp      (io_node_axi_1_b_payload_resp[1:0]         ), //i
    .io_axi_1_ar_valid            (nodeFlow_io_axi_1_ar_valid                ), //o
    .io_axi_1_ar_ready            (io_node_axi_1_ar_ready                    ), //i
    .io_axi_1_ar_payload_addr     (nodeFlow_io_axi_1_ar_payload_addr[63:0]   ), //o
    .io_axi_1_ar_payload_id       (nodeFlow_io_axi_1_ar_payload_id[5:0]      ), //o
    .io_axi_1_ar_payload_len      (nodeFlow_io_axi_1_ar_payload_len[7:0]     ), //o
    .io_axi_1_ar_payload_size     (nodeFlow_io_axi_1_ar_payload_size[2:0]    ), //o
    .io_axi_1_ar_payload_burst    (nodeFlow_io_axi_1_ar_payload_burst[1:0]   ), //o
    .io_axi_1_r_valid             (io_node_axi_1_r_valid                     ), //i
    .io_axi_1_r_ready             (nodeFlow_io_axi_1_r_ready                 ), //o
    .io_axi_1_r_payload_data      (io_node_axi_1_r_payload_data[511:0]       ), //i
    .io_axi_1_r_payload_id        (io_node_axi_1_r_payload_id[5:0]           ), //i
    .io_axi_1_r_payload_resp      (io_node_axi_1_r_payload_resp[1:0]         ), //i
    .io_axi_1_r_payload_last      (io_node_axi_1_r_payload_last              ), //i
    .io_cmdAxi_0_aw_valid         (nodeFlow_io_cmdAxi_0_aw_valid             ), //o
    .io_cmdAxi_0_aw_ready         (io_node_cmdAxi_0_aw_ready                 ), //i
    .io_cmdAxi_0_aw_payload_addr  (nodeFlow_io_cmdAxi_0_aw_payload_addr[63:0]), //o
    .io_cmdAxi_0_aw_payload_id    (nodeFlow_io_cmdAxi_0_aw_payload_id[5:0]   ), //o
    .io_cmdAxi_0_aw_payload_len   (nodeFlow_io_cmdAxi_0_aw_payload_len[7:0]  ), //o
    .io_cmdAxi_0_aw_payload_size  (nodeFlow_io_cmdAxi_0_aw_payload_size[2:0] ), //o
    .io_cmdAxi_0_aw_payload_burst (nodeFlow_io_cmdAxi_0_aw_payload_burst[1:0]), //o
    .io_cmdAxi_0_w_valid          (nodeFlow_io_cmdAxi_0_w_valid              ), //o
    .io_cmdAxi_0_w_ready          (io_node_cmdAxi_0_w_ready                  ), //i
    .io_cmdAxi_0_w_payload_data   (nodeFlow_io_cmdAxi_0_w_payload_data[511:0]), //o
    .io_cmdAxi_0_w_payload_strb   (nodeFlow_io_cmdAxi_0_w_payload_strb[63:0] ), //o
    .io_cmdAxi_0_w_payload_last   (nodeFlow_io_cmdAxi_0_w_payload_last       ), //o
    .io_cmdAxi_0_b_valid          (io_node_cmdAxi_0_b_valid                  ), //i
    .io_cmdAxi_0_b_ready          (nodeFlow_io_cmdAxi_0_b_ready              ), //o
    .io_cmdAxi_0_b_payload_id     (io_node_cmdAxi_0_b_payload_id[5:0]        ), //i
    .io_cmdAxi_0_b_payload_resp   (io_node_cmdAxi_0_b_payload_resp[1:0]      ), //i
    .io_cmdAxi_0_ar_valid         (nodeFlow_io_cmdAxi_0_ar_valid             ), //o
    .io_cmdAxi_0_ar_ready         (io_node_cmdAxi_0_ar_ready                 ), //i
    .io_cmdAxi_0_ar_payload_addr  (nodeFlow_io_cmdAxi_0_ar_payload_addr[63:0]), //o
    .io_cmdAxi_0_ar_payload_id    (nodeFlow_io_cmdAxi_0_ar_payload_id[5:0]   ), //o
    .io_cmdAxi_0_ar_payload_len   (nodeFlow_io_cmdAxi_0_ar_payload_len[7:0]  ), //o
    .io_cmdAxi_0_ar_payload_size  (nodeFlow_io_cmdAxi_0_ar_payload_size[2:0] ), //o
    .io_cmdAxi_0_ar_payload_burst (nodeFlow_io_cmdAxi_0_ar_payload_burst[1:0]), //o
    .io_cmdAxi_0_r_valid          (io_node_cmdAxi_0_r_valid                  ), //i
    .io_cmdAxi_0_r_ready          (nodeFlow_io_cmdAxi_0_r_ready              ), //o
    .io_cmdAxi_0_r_payload_data   (io_node_cmdAxi_0_r_payload_data[511:0]    ), //i
    .io_cmdAxi_0_r_payload_id     (io_node_cmdAxi_0_r_payload_id[5:0]        ), //i
    .io_cmdAxi_0_r_payload_resp   (io_node_cmdAxi_0_r_payload_resp[1:0]      ), //i
    .io_cmdAxi_0_r_payload_last   (io_node_cmdAxi_0_r_payload_last           ), //i
    .io_nodeId                    (io_node_nodeId                            ), //i
    .io_txnNumTotal               (io_node_txnNumTotal[31:0]                 ), //i
    .io_cmdAddrOffs_0             (io_node_cmdAddrOffs_0[31:0]               ), //i
    .io_start                     (io_node_start                             ), //i
    .io_done_0                    (nodeFlow_io_done_0                        ), //o
    .io_cntTxnCmt_0               (nodeFlow_io_cntTxnCmt_0[31:0]             ), //o
    .io_cntTxnAbt_0               (nodeFlow_io_cntTxnAbt_0[31:0]             ), //o
    .io_cntTxnLd_0                (nodeFlow_io_cntTxnLd_0[31:0]              ), //o
    .io_cntLockLoc_0              (nodeFlow_io_cntLockLoc_0[31:0]            ), //o
    .io_cntLockRmt_0              (nodeFlow_io_cntLockRmt_0[31:0]            ), //o
    .io_cntLockDenyLoc_0          (nodeFlow_io_cntLockDenyLoc_0[31:0]        ), //o
    .io_cntLockDenyRmt_0          (nodeFlow_io_cntLockDenyRmt_0[31:0]        ), //o
    .io_cntClk_0                  (nodeFlow_io_cntClk_0[31:0]                ), //o
    .io_sendQ_valid               (nodeFlow_io_sendQ_valid                   ), //o
    .io_sendQ_ready               (rdmaFlowMstr_io_q_sink_ready              ), //i
    .io_sendQ_payload             (nodeFlow_io_sendQ_payload[511:0]          ), //o
    .io_respQ_valid               (nodeFlow_io_respQ_valid                   ), //o
    .io_respQ_ready               (rdmaFlowSlve_io_q_sink_ready              ), //i
    .io_respQ_payload             (nodeFlow_io_respQ_payload[511:0]          ), //o
    .io_reqQ_valid                (rdmaFlowSlve_io_q_src_valid               ), //i
    .io_reqQ_ready                (nodeFlow_io_reqQ_ready                    ), //o
    .io_reqQ_payload              (rdmaFlowSlve_io_q_src_payload[511:0]      ), //i
    .io_recvQ_valid               (rdmaFlowMstr_io_q_src_valid               ), //i
    .io_recvQ_ready               (nodeFlow_io_recvQ_ready                   ), //o
    .io_recvQ_payload             (rdmaFlowMstr_io_q_src_payload[511:0]      ), //i
    .io_sendStatusVld             (nodeFlow_io_sendStatusVld                 ), //o
    .io_recvStatusVld             (nodeFlow_io_recvStatusVld                 ), //o
    .io_nReq                      (nodeFlow_io_nReq[3:0]                     ), //o
    .io_nWrCmtReq                 (nodeFlow_io_nWrCmtReq[3:0]                ), //o
    .io_nRdGetReq                 (nodeFlow_io_nRdGetReq[3:0]                ), //o
    .io_nResp                     (nodeFlow_io_nResp[3:0]                    ), //o
    .io_nWrCmtResp                (nodeFlow_io_nWrCmtResp[3:0]               ), //o
    .io_nRdGetResp                (nodeFlow_io_nRdGetResp[3:0]               ), //o
    .resetn                       (resetn                                    ), //i
    .clk                          (clk                                       )  //i
  );
  RdmaFlowBpss rdmaFlowMstr (
    .io_rdma_rd_req_valid            (rdmaArb_1_io_rdmaV_0_rd_req_valid                  ), //i
    .io_rdma_rd_req_ready            (rdmaFlowMstr_io_rdma_rd_req_ready                  ), //o
    .io_rdma_rd_req_payload_data     (rdmaArb_1_io_rdmaV_0_rd_req_payload_data[95:0]     ), //i
    .io_rdma_wr_req_valid            (rdmaArb_1_io_rdmaV_0_wr_req_valid                  ), //i
    .io_rdma_wr_req_ready            (rdmaFlowMstr_io_rdma_wr_req_ready                  ), //o
    .io_rdma_wr_req_payload_data     (rdmaArb_1_io_rdmaV_0_wr_req_payload_data[95:0]     ), //i
    .io_rdma_sq_valid                (rdmaFlowMstr_io_rdma_sq_valid                      ), //o
    .io_rdma_sq_ready                (rdmaArb_1_io_rdmaV_0_sq_ready                      ), //i
    .io_rdma_sq_payload_data         (rdmaFlowMstr_io_rdma_sq_payload_data[543:0]        ), //o
    .io_rdma_ack_valid               (rdmaArb_1_io_rdmaV_0_ack_valid                     ), //i
    .io_rdma_ack_ready               (rdmaFlowMstr_io_rdma_ack_ready                     ), //o
    .io_rdma_ack_payload_data        (rdmaArb_1_io_rdmaV_0_ack_payload_data[42:0]        ), //i
    .io_rdma_axis_sink_valid         (rdmaArb_1_io_rdmaV_0_axis_sink_valid               ), //i
    .io_rdma_axis_sink_ready         (rdmaFlowMstr_io_rdma_axis_sink_ready               ), //o
    .io_rdma_axis_sink_payload_tdata (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tdata[511:0]), //i
    .io_rdma_axis_sink_payload_tkeep (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tkeep[63:0] ), //i
    .io_rdma_axis_sink_payload_tlast (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tlast       ), //i
    .io_rdma_axis_src_valid          (rdmaFlowMstr_io_rdma_axis_src_valid                ), //o
    .io_rdma_axis_src_ready          (rdmaArb_1_io_rdmaV_0_axis_src_ready                ), //i
    .io_rdma_axis_src_payload_tdata  (rdmaFlowMstr_io_rdma_axis_src_payload_tdata[511:0] ), //o
    .io_rdma_axis_src_payload_tkeep  (rdmaFlowMstr_io_rdma_axis_src_payload_tkeep[63:0]  ), //o
    .io_rdma_axis_src_payload_tlast  (rdmaFlowMstr_io_rdma_axis_src_payload_tlast        ), //o
    .io_q_sink_valid                 (nodeFlow_io_sendQ_valid                            ), //i
    .io_q_sink_ready                 (rdmaFlowMstr_io_q_sink_ready                       ), //o
    .io_q_sink_payload               (nodeFlow_io_sendQ_payload[511:0]                   ), //i
    .io_q_src_valid                  (rdmaFlowMstr_io_q_src_valid                        ), //o
    .io_q_src_ready                  (nodeFlow_io_recvQ_ready                            ), //i
    .io_q_src_payload                (rdmaFlowMstr_io_q_src_payload[511:0]               ), //o
    .io_ctrl_en                      (io_rdmaCtrl_0_en                                   ), //i
    .io_ctrl_len                     (io_rdmaCtrl_0_len[31:0]                            ), //i
    .io_ctrl_qpn                     (io_rdmaCtrl_0_qpn[9:0]                             ), //i
    .io_ctrl_flowId                  (io_rdmaCtrl_0_flowId[3:0]                          ), //i
    .clk                             (clk                                                ), //i
    .resetn                          (resetn                                             )  //i
  );
  RdmaFlowBpss_1 rdmaFlowSlve (
    .io_rdma_rd_req_valid            (rdmaArb_1_io_rdmaV_1_rd_req_valid                  ), //i
    .io_rdma_rd_req_ready            (rdmaFlowSlve_io_rdma_rd_req_ready                  ), //o
    .io_rdma_rd_req_payload_data     (rdmaArb_1_io_rdmaV_1_rd_req_payload_data[95:0]     ), //i
    .io_rdma_wr_req_valid            (rdmaArb_1_io_rdmaV_1_wr_req_valid                  ), //i
    .io_rdma_wr_req_ready            (rdmaFlowSlve_io_rdma_wr_req_ready                  ), //o
    .io_rdma_wr_req_payload_data     (rdmaArb_1_io_rdmaV_1_wr_req_payload_data[95:0]     ), //i
    .io_rdma_sq_valid                (rdmaFlowSlve_io_rdma_sq_valid                      ), //o
    .io_rdma_sq_ready                (rdmaArb_1_io_rdmaV_1_sq_ready                      ), //i
    .io_rdma_sq_payload_data         (rdmaFlowSlve_io_rdma_sq_payload_data[543:0]        ), //o
    .io_rdma_ack_valid               (rdmaArb_1_io_rdmaV_1_ack_valid                     ), //i
    .io_rdma_ack_ready               (rdmaFlowSlve_io_rdma_ack_ready                     ), //o
    .io_rdma_ack_payload_data        (rdmaArb_1_io_rdmaV_1_ack_payload_data[42:0]        ), //i
    .io_rdma_axis_sink_valid         (rdmaArb_1_io_rdmaV_1_axis_sink_valid               ), //i
    .io_rdma_axis_sink_ready         (rdmaFlowSlve_io_rdma_axis_sink_ready               ), //o
    .io_rdma_axis_sink_payload_tdata (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tdata[511:0]), //i
    .io_rdma_axis_sink_payload_tkeep (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tkeep[63:0] ), //i
    .io_rdma_axis_sink_payload_tlast (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tlast       ), //i
    .io_rdma_axis_src_valid          (rdmaFlowSlve_io_rdma_axis_src_valid                ), //o
    .io_rdma_axis_src_ready          (rdmaArb_1_io_rdmaV_1_axis_src_ready                ), //i
    .io_rdma_axis_src_payload_tdata  (rdmaFlowSlve_io_rdma_axis_src_payload_tdata[511:0] ), //o
    .io_rdma_axis_src_payload_tkeep  (rdmaFlowSlve_io_rdma_axis_src_payload_tkeep[63:0]  ), //o
    .io_rdma_axis_src_payload_tlast  (rdmaFlowSlve_io_rdma_axis_src_payload_tlast        ), //o
    .io_q_sink_valid                 (nodeFlow_io_respQ_valid                            ), //i
    .io_q_sink_ready                 (rdmaFlowSlve_io_q_sink_ready                       ), //o
    .io_q_sink_payload               (nodeFlow_io_respQ_payload[511:0]                   ), //i
    .io_q_src_valid                  (rdmaFlowSlve_io_q_src_valid                        ), //o
    .io_q_src_ready                  (nodeFlow_io_reqQ_ready                             ), //i
    .io_q_src_payload                (rdmaFlowSlve_io_q_src_payload[511:0]               ), //o
    .io_ctrl_en                      (io_rdmaCtrl_1_en                                   ), //i
    .io_ctrl_len                     (io_rdmaCtrl_1_len[31:0]                            ), //i
    .io_ctrl_qpn                     (io_rdmaCtrl_1_qpn[9:0]                             ), //i
    .io_ctrl_flowId                  (io_rdmaCtrl_1_flowId[3:0]                          ), //i
    .clk                             (clk                                                ), //i
    .resetn                          (resetn                                             )  //i
  );
  RdmaArb rdmaArb_1 (
    .io_rdmaV_0_rd_req_valid            (rdmaArb_1_io_rdmaV_0_rd_req_valid                  ), //o
    .io_rdmaV_0_rd_req_ready            (rdmaFlowMstr_io_rdma_rd_req_ready                  ), //i
    .io_rdmaV_0_rd_req_payload_data     (rdmaArb_1_io_rdmaV_0_rd_req_payload_data[95:0]     ), //o
    .io_rdmaV_0_wr_req_valid            (rdmaArb_1_io_rdmaV_0_wr_req_valid                  ), //o
    .io_rdmaV_0_wr_req_ready            (rdmaFlowMstr_io_rdma_wr_req_ready                  ), //i
    .io_rdmaV_0_wr_req_payload_data     (rdmaArb_1_io_rdmaV_0_wr_req_payload_data[95:0]     ), //o
    .io_rdmaV_0_sq_valid                (rdmaFlowMstr_io_rdma_sq_valid                      ), //i
    .io_rdmaV_0_sq_ready                (rdmaArb_1_io_rdmaV_0_sq_ready                      ), //o
    .io_rdmaV_0_sq_payload_data         (rdmaFlowMstr_io_rdma_sq_payload_data[543:0]        ), //i
    .io_rdmaV_0_ack_valid               (rdmaArb_1_io_rdmaV_0_ack_valid                     ), //o
    .io_rdmaV_0_ack_ready               (rdmaFlowMstr_io_rdma_ack_ready                     ), //i
    .io_rdmaV_0_ack_payload_data        (rdmaArb_1_io_rdmaV_0_ack_payload_data[42:0]        ), //o
    .io_rdmaV_0_axis_sink_valid         (rdmaArb_1_io_rdmaV_0_axis_sink_valid               ), //o
    .io_rdmaV_0_axis_sink_ready         (rdmaFlowMstr_io_rdma_axis_sink_ready               ), //i
    .io_rdmaV_0_axis_sink_payload_tdata (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tdata[511:0]), //o
    .io_rdmaV_0_axis_sink_payload_tkeep (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tkeep[63:0] ), //o
    .io_rdmaV_0_axis_sink_payload_tlast (rdmaArb_1_io_rdmaV_0_axis_sink_payload_tlast       ), //o
    .io_rdmaV_0_axis_src_valid          (rdmaFlowMstr_io_rdma_axis_src_valid                ), //i
    .io_rdmaV_0_axis_src_ready          (rdmaArb_1_io_rdmaV_0_axis_src_ready                ), //o
    .io_rdmaV_0_axis_src_payload_tdata  (rdmaFlowMstr_io_rdma_axis_src_payload_tdata[511:0] ), //i
    .io_rdmaV_0_axis_src_payload_tkeep  (rdmaFlowMstr_io_rdma_axis_src_payload_tkeep[63:0]  ), //i
    .io_rdmaV_0_axis_src_payload_tlast  (rdmaFlowMstr_io_rdma_axis_src_payload_tlast        ), //i
    .io_rdmaV_1_rd_req_valid            (rdmaArb_1_io_rdmaV_1_rd_req_valid                  ), //o
    .io_rdmaV_1_rd_req_ready            (rdmaFlowSlve_io_rdma_rd_req_ready                  ), //i
    .io_rdmaV_1_rd_req_payload_data     (rdmaArb_1_io_rdmaV_1_rd_req_payload_data[95:0]     ), //o
    .io_rdmaV_1_wr_req_valid            (rdmaArb_1_io_rdmaV_1_wr_req_valid                  ), //o
    .io_rdmaV_1_wr_req_ready            (rdmaFlowSlve_io_rdma_wr_req_ready                  ), //i
    .io_rdmaV_1_wr_req_payload_data     (rdmaArb_1_io_rdmaV_1_wr_req_payload_data[95:0]     ), //o
    .io_rdmaV_1_sq_valid                (rdmaFlowSlve_io_rdma_sq_valid                      ), //i
    .io_rdmaV_1_sq_ready                (rdmaArb_1_io_rdmaV_1_sq_ready                      ), //o
    .io_rdmaV_1_sq_payload_data         (rdmaFlowSlve_io_rdma_sq_payload_data[543:0]        ), //i
    .io_rdmaV_1_ack_valid               (rdmaArb_1_io_rdmaV_1_ack_valid                     ), //o
    .io_rdmaV_1_ack_ready               (rdmaFlowSlve_io_rdma_ack_ready                     ), //i
    .io_rdmaV_1_ack_payload_data        (rdmaArb_1_io_rdmaV_1_ack_payload_data[42:0]        ), //o
    .io_rdmaV_1_axis_sink_valid         (rdmaArb_1_io_rdmaV_1_axis_sink_valid               ), //o
    .io_rdmaV_1_axis_sink_ready         (rdmaFlowSlve_io_rdma_axis_sink_ready               ), //i
    .io_rdmaV_1_axis_sink_payload_tdata (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tdata[511:0]), //o
    .io_rdmaV_1_axis_sink_payload_tkeep (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tkeep[63:0] ), //o
    .io_rdmaV_1_axis_sink_payload_tlast (rdmaArb_1_io_rdmaV_1_axis_sink_payload_tlast       ), //o
    .io_rdmaV_1_axis_src_valid          (rdmaFlowSlve_io_rdma_axis_src_valid                ), //i
    .io_rdmaV_1_axis_src_ready          (rdmaArb_1_io_rdmaV_1_axis_src_ready                ), //o
    .io_rdmaV_1_axis_src_payload_tdata  (rdmaFlowSlve_io_rdma_axis_src_payload_tdata[511:0] ), //i
    .io_rdmaV_1_axis_src_payload_tkeep  (rdmaFlowSlve_io_rdma_axis_src_payload_tkeep[63:0]  ), //i
    .io_rdmaV_1_axis_src_payload_tlast  (rdmaFlowSlve_io_rdma_axis_src_payload_tlast        ), //i
    .io_rdmaio_rd_req_valid             (io_rdma_rd_req_valid                               ), //i
    .io_rdmaio_rd_req_ready             (rdmaArb_1_io_rdmaio_rd_req_ready                   ), //o
    .io_rdmaio_rd_req_payload_data      (io_rdma_rd_req_payload_data[95:0]                  ), //i
    .io_rdmaio_wr_req_valid             (io_rdma_wr_req_valid                               ), //i
    .io_rdmaio_wr_req_ready             (rdmaArb_1_io_rdmaio_wr_req_ready                   ), //o
    .io_rdmaio_wr_req_payload_data      (io_rdma_wr_req_payload_data[95:0]                  ), //i
    .io_rdmaio_sq_valid                 (rdmaArb_1_io_rdmaio_sq_valid                       ), //o
    .io_rdmaio_sq_ready                 (io_rdma_sq_ready                                   ), //i
    .io_rdmaio_sq_payload_data          (rdmaArb_1_io_rdmaio_sq_payload_data[543:0]         ), //o
    .io_rdmaio_ack_valid                (io_rdma_ack_valid                                  ), //i
    .io_rdmaio_ack_ready                (rdmaArb_1_io_rdmaio_ack_ready                      ), //o
    .io_rdmaio_ack_payload_data         (io_rdma_ack_payload_data[42:0]                     ), //i
    .io_rdmaio_axis_sink_valid          (io_rdma_axis_sink_valid                            ), //i
    .io_rdmaio_axis_sink_ready          (rdmaArb_1_io_rdmaio_axis_sink_ready                ), //o
    .io_rdmaio_axis_sink_payload_tdata  (io_rdma_axis_sink_payload_tdata[511:0]             ), //i
    .io_rdmaio_axis_sink_payload_tkeep  (io_rdma_axis_sink_payload_tkeep[63:0]              ), //i
    .io_rdmaio_axis_sink_payload_tlast  (io_rdma_axis_sink_payload_tlast                    ), //i
    .io_rdmaio_axis_src_valid           (rdmaArb_1_io_rdmaio_axis_src_valid                 ), //o
    .io_rdmaio_axis_src_ready           (io_rdma_axis_src_ready                             ), //i
    .io_rdmaio_axis_src_payload_tdata   (rdmaArb_1_io_rdmaio_axis_src_payload_tdata[511:0]  ), //o
    .io_rdmaio_axis_src_payload_tkeep   (rdmaArb_1_io_rdmaio_axis_src_payload_tkeep[63:0]   ), //o
    .io_rdmaio_axis_src_payload_tlast   (rdmaArb_1_io_rdmaio_axis_src_payload_tlast         ), //o
    .clk                                (clk                                                ), //i
    .resetn                             (resetn                                             )  //i
  );
  assign io_node_axi_0_aw_valid = nodeFlow_io_axi_0_aw_valid;
  assign io_node_axi_0_aw_payload_addr = nodeFlow_io_axi_0_aw_payload_addr;
  assign io_node_axi_0_aw_payload_id = nodeFlow_io_axi_0_aw_payload_id;
  assign io_node_axi_0_aw_payload_len = nodeFlow_io_axi_0_aw_payload_len;
  assign io_node_axi_0_aw_payload_size = nodeFlow_io_axi_0_aw_payload_size;
  assign io_node_axi_0_aw_payload_burst = nodeFlow_io_axi_0_aw_payload_burst;
  assign io_node_axi_0_w_valid = nodeFlow_io_axi_0_w_valid;
  assign io_node_axi_0_w_payload_data = nodeFlow_io_axi_0_w_payload_data;
  assign io_node_axi_0_w_payload_strb = nodeFlow_io_axi_0_w_payload_strb;
  assign io_node_axi_0_w_payload_last = nodeFlow_io_axi_0_w_payload_last;
  assign io_node_axi_0_b_ready = nodeFlow_io_axi_0_b_ready;
  assign io_node_axi_0_ar_valid = nodeFlow_io_axi_0_ar_valid;
  assign io_node_axi_0_ar_payload_addr = nodeFlow_io_axi_0_ar_payload_addr;
  assign io_node_axi_0_ar_payload_id = nodeFlow_io_axi_0_ar_payload_id;
  assign io_node_axi_0_ar_payload_len = nodeFlow_io_axi_0_ar_payload_len;
  assign io_node_axi_0_ar_payload_size = nodeFlow_io_axi_0_ar_payload_size;
  assign io_node_axi_0_ar_payload_burst = nodeFlow_io_axi_0_ar_payload_burst;
  assign io_node_axi_0_r_ready = nodeFlow_io_axi_0_r_ready;
  assign io_node_axi_1_aw_valid = nodeFlow_io_axi_1_aw_valid;
  assign io_node_axi_1_aw_payload_addr = nodeFlow_io_axi_1_aw_payload_addr;
  assign io_node_axi_1_aw_payload_id = nodeFlow_io_axi_1_aw_payload_id;
  assign io_node_axi_1_aw_payload_len = nodeFlow_io_axi_1_aw_payload_len;
  assign io_node_axi_1_aw_payload_size = nodeFlow_io_axi_1_aw_payload_size;
  assign io_node_axi_1_aw_payload_burst = nodeFlow_io_axi_1_aw_payload_burst;
  assign io_node_axi_1_w_valid = nodeFlow_io_axi_1_w_valid;
  assign io_node_axi_1_w_payload_data = nodeFlow_io_axi_1_w_payload_data;
  assign io_node_axi_1_w_payload_strb = nodeFlow_io_axi_1_w_payload_strb;
  assign io_node_axi_1_w_payload_last = nodeFlow_io_axi_1_w_payload_last;
  assign io_node_axi_1_b_ready = nodeFlow_io_axi_1_b_ready;
  assign io_node_axi_1_ar_valid = nodeFlow_io_axi_1_ar_valid;
  assign io_node_axi_1_ar_payload_addr = nodeFlow_io_axi_1_ar_payload_addr;
  assign io_node_axi_1_ar_payload_id = nodeFlow_io_axi_1_ar_payload_id;
  assign io_node_axi_1_ar_payload_len = nodeFlow_io_axi_1_ar_payload_len;
  assign io_node_axi_1_ar_payload_size = nodeFlow_io_axi_1_ar_payload_size;
  assign io_node_axi_1_ar_payload_burst = nodeFlow_io_axi_1_ar_payload_burst;
  assign io_node_axi_1_r_ready = nodeFlow_io_axi_1_r_ready;
  assign io_node_cmdAxi_0_aw_valid = nodeFlow_io_cmdAxi_0_aw_valid;
  assign io_node_cmdAxi_0_aw_payload_addr = nodeFlow_io_cmdAxi_0_aw_payload_addr;
  assign io_node_cmdAxi_0_aw_payload_id = nodeFlow_io_cmdAxi_0_aw_payload_id;
  assign io_node_cmdAxi_0_aw_payload_len = nodeFlow_io_cmdAxi_0_aw_payload_len;
  assign io_node_cmdAxi_0_aw_payload_size = nodeFlow_io_cmdAxi_0_aw_payload_size;
  assign io_node_cmdAxi_0_aw_payload_burst = nodeFlow_io_cmdAxi_0_aw_payload_burst;
  assign io_node_cmdAxi_0_w_valid = nodeFlow_io_cmdAxi_0_w_valid;
  assign io_node_cmdAxi_0_w_payload_data = nodeFlow_io_cmdAxi_0_w_payload_data;
  assign io_node_cmdAxi_0_w_payload_strb = nodeFlow_io_cmdAxi_0_w_payload_strb;
  assign io_node_cmdAxi_0_w_payload_last = nodeFlow_io_cmdAxi_0_w_payload_last;
  assign io_node_cmdAxi_0_b_ready = nodeFlow_io_cmdAxi_0_b_ready;
  assign io_node_cmdAxi_0_ar_valid = nodeFlow_io_cmdAxi_0_ar_valid;
  assign io_node_cmdAxi_0_ar_payload_addr = nodeFlow_io_cmdAxi_0_ar_payload_addr;
  assign io_node_cmdAxi_0_ar_payload_id = nodeFlow_io_cmdAxi_0_ar_payload_id;
  assign io_node_cmdAxi_0_ar_payload_len = nodeFlow_io_cmdAxi_0_ar_payload_len;
  assign io_node_cmdAxi_0_ar_payload_size = nodeFlow_io_cmdAxi_0_ar_payload_size;
  assign io_node_cmdAxi_0_ar_payload_burst = nodeFlow_io_cmdAxi_0_ar_payload_burst;
  assign io_node_cmdAxi_0_r_ready = nodeFlow_io_cmdAxi_0_r_ready;
  assign io_node_done_0 = nodeFlow_io_done_0;
  assign io_node_cntTxnCmt_0 = nodeFlow_io_cntTxnCmt_0;
  assign io_node_cntTxnAbt_0 = nodeFlow_io_cntTxnAbt_0;
  assign io_node_cntTxnLd_0 = nodeFlow_io_cntTxnLd_0;
  assign io_node_cntLockLoc_0 = nodeFlow_io_cntLockLoc_0;
  assign io_node_cntLockRmt_0 = nodeFlow_io_cntLockRmt_0;
  assign io_node_cntLockDenyLoc_0 = nodeFlow_io_cntLockDenyLoc_0;
  assign io_node_cntLockDenyRmt_0 = nodeFlow_io_cntLockDenyRmt_0;
  assign io_node_cntClk_0 = nodeFlow_io_cntClk_0;
  assign io_rdma_rd_req_ready = rdmaArb_1_io_rdmaio_rd_req_ready;
  assign io_rdma_wr_req_ready = rdmaArb_1_io_rdmaio_wr_req_ready;
  assign io_rdma_sq_valid = rdmaArb_1_io_rdmaio_sq_valid;
  assign io_rdma_sq_payload_data = rdmaArb_1_io_rdmaio_sq_payload_data;
  assign io_rdma_ack_ready = rdmaArb_1_io_rdmaio_ack_ready;
  assign io_rdma_axis_sink_ready = rdmaArb_1_io_rdmaio_axis_sink_ready;
  assign io_rdma_axis_src_valid = rdmaArb_1_io_rdmaio_axis_src_valid;
  assign io_rdma_axis_src_payload_tdata = rdmaArb_1_io_rdmaio_axis_src_payload_tdata;
  assign io_rdma_axis_src_payload_tkeep = rdmaArb_1_io_rdmaio_axis_src_payload_tkeep;
  assign io_rdma_axis_src_payload_tlast = rdmaArb_1_io_rdmaio_axis_src_payload_tlast;
  always @(*) begin
    cntSent_willIncrement = 1'b0;
    if(io_rdma_axis_src_fire) begin
      cntSent_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    cntSent_willClear = 1'b0;
    if(when_WrapNodeNet_l49) begin
      cntSent_willClear = 1'b1;
    end
  end

  assign cntSent_willOverflowIfInc = (cntSent_value == 32'hffffffff);
  assign cntSent_willOverflow = (cntSent_willOverflowIfInc && cntSent_willIncrement);
  always @(*) begin
    cntSent_valueNext = (cntSent_value + _zz_cntSent_valueNext);
    if(cntSent_willClear) begin
      cntSent_valueNext = 32'h0;
    end
  end

  always @(*) begin
    cntRecv_willIncrement = 1'b0;
    if(io_rdma_axis_sink_fire) begin
      cntRecv_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    cntRecv_willClear = 1'b0;
    if(when_WrapNodeNet_l52) begin
      cntRecv_willClear = 1'b1;
    end
  end

  assign cntRecv_willOverflowIfInc = (cntRecv_value == 32'hffffffff);
  assign cntRecv_willOverflow = (cntRecv_willOverflowIfInc && cntRecv_willIncrement);
  always @(*) begin
    cntRecv_valueNext = (cntRecv_value + _zz_cntRecv_valueNext);
    if(cntRecv_willClear) begin
      cntRecv_valueNext = 32'h0;
    end
  end

  assign io_rdma_axis_src_fire = (io_rdma_axis_src_valid && io_rdma_axis_src_ready);
  assign io_rdma_axis_sink_fire = (io_rdma_axis_sink_valid && io_rdma_axis_sink_ready);
  assign when_WrapNodeNet_l49 = (! io_rdmaCtrl_0_en);
  assign when_WrapNodeNet_l52 = (! io_rdmaCtrl_1_en);
  assign io_cntRDMASent = cntSent_value;
  assign io_cntRDMARecv = cntRecv_value;
  always @(posedge clk) begin
    if(!resetn) begin
      cntSent_value <= 32'h0;
      cntRecv_value <= 32'h0;
    end else begin
      cntSent_value <= cntSent_valueNext;
      cntRecv_value <= cntRecv_valueNext;
    end
  end


endmodule

module CMemHost (
  input      [1:0]    io_mode,
  input      [63:0]   io_hostAddr,
  input      [63:0]   io_cmemAddr,
  input      [15:0]   io_len,
  input      [63:0]   io_cnt,
  input      [5:0]    io_pid,
  output reg [63:0]   io_cntDone,
  output              io_hostd_bpss_rd_req_valid,
  input               io_hostd_bpss_rd_req_ready,
  output     [95:0]   io_hostd_bpss_rd_req_payload_data,
  output              io_hostd_bpss_wr_req_valid,
  input               io_hostd_bpss_wr_req_ready,
  output     [95:0]   io_hostd_bpss_wr_req_payload_data,
  input               io_hostd_bpss_rd_done_valid,
  output              io_hostd_bpss_rd_done_ready,
  input      [5:0]    io_hostd_bpss_rd_done_payload_data,
  input               io_hostd_bpss_wr_done_valid,
  output              io_hostd_bpss_wr_done_ready,
  input      [5:0]    io_hostd_bpss_wr_done_payload_data,
  input               io_hostd_axis_host_sink_valid,
  output              io_hostd_axis_host_sink_ready,
  input      [511:0]  io_hostd_axis_host_sink_payload_tdata,
  input      [3:0]    io_hostd_axis_host_sink_payload_tdest,
  input      [63:0]   io_hostd_axis_host_sink_payload_tkeep,
  input               io_hostd_axis_host_sink_payload_tlast,
  output              io_hostd_axis_host_src_valid,
  input               io_hostd_axis_host_src_ready,
  output     [511:0]  io_hostd_axis_host_src_payload_tdata,
  output     [3:0]    io_hostd_axis_host_src_payload_tdest,
  output     [63:0]   io_hostd_axis_host_src_payload_tkeep,
  output              io_hostd_axis_host_src_payload_tlast,
  output              io_axi_cmem_aw_valid,
  input               io_axi_cmem_aw_ready,
  output     [63:0]   io_axi_cmem_aw_payload_addr,
  output     [5:0]    io_axi_cmem_aw_payload_id,
  output     [7:0]    io_axi_cmem_aw_payload_len,
  output     [2:0]    io_axi_cmem_aw_payload_size,
  output     [1:0]    io_axi_cmem_aw_payload_burst,
  output              io_axi_cmem_w_valid,
  input               io_axi_cmem_w_ready,
  output     [511:0]  io_axi_cmem_w_payload_data,
  output     [63:0]   io_axi_cmem_w_payload_strb,
  output              io_axi_cmem_w_payload_last,
  input               io_axi_cmem_b_valid,
  output              io_axi_cmem_b_ready,
  input      [5:0]    io_axi_cmem_b_payload_id,
  input      [1:0]    io_axi_cmem_b_payload_resp,
  output              io_axi_cmem_ar_valid,
  input               io_axi_cmem_ar_ready,
  output     [63:0]   io_axi_cmem_ar_payload_addr,
  output     [5:0]    io_axi_cmem_ar_payload_id,
  output     [7:0]    io_axi_cmem_ar_payload_len,
  output     [2:0]    io_axi_cmem_ar_payload_size,
  output     [1:0]    io_axi_cmem_ar_payload_burst,
  input               io_axi_cmem_r_valid,
  output              io_axi_cmem_r_ready,
  input      [511:0]  io_axi_cmem_r_payload_data,
  input      [5:0]    io_axi_cmem_r_payload_id,
  input      [1:0]    io_axi_cmem_r_payload_resp,
  input               io_axi_cmem_r_payload_last,
  input               clk,
  input               resetn
);
  localparam fsm_enumDef_BOOT = 2'd0;
  localparam fsm_enumDef_IDLE = 2'd1;
  localparam fsm_enumDef_RD = 2'd2;
  localparam fsm_enumDef_WR = 2'd3;

  wire       [63:0]   _zz_reqHostAddr;
  wire       [9:0]    _zz_io_axi_cmem_aw_payload_len;
  wire       [9:0]    _zz_io_axi_cmem_aw_payload_len_1;
  wire       [9:0]    _zz_io_axi_cmem_ar_payload_len;
  wire       [9:0]    _zz_io_axi_cmem_ar_payload_len_1;
  wire       [63:0]   _zz_cmemWrAddr;
  wire       [63:0]   _zz_cmemRdAddr;
  reg        [63:0]   cntWrData;
  reg        [63:0]   cntRdData;
  reg        [63:0]   cntHostReq;
  reg        [63:0]   cntHbmReq;
  reg        [63:0]   cmemRdAddr;
  reg        [63:0]   cmemWrAddr;
  reg        [63:0]   reqHostAddr;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  wire       [4:0]    bpss_rd_req_rsrvd;
  wire       [0:0]    bpss_rd_req_vfid;
  wire       [5:0]    bpss_rd_req_pid;
  wire       [3:0]    bpss_rd_req_dest;
  wire                bpss_rd_req_host;
  wire                bpss_rd_req_ctl;
  wire                bpss_rd_req_sync;
  wire                bpss_rd_req_stream;
  wire       [27:0]   bpss_rd_req_len;
  wire       [47:0]   bpss_rd_req_vaddr;
  wire       [4:0]    bpss_wr_req_rsrvd;
  wire       [0:0]    bpss_wr_req_vfid;
  wire       [5:0]    bpss_wr_req_pid;
  wire       [3:0]    bpss_wr_req_dest;
  wire                bpss_wr_req_host;
  wire                bpss_wr_req_ctl;
  wire                bpss_wr_req_sync;
  wire                bpss_wr_req_stream;
  wire       [27:0]   bpss_wr_req_len;
  wire       [47:0]   bpss_wr_req_vaddr;
  wire                io_hostd_bpss_rd_req_fire;
  wire                io_hostd_bpss_wr_req_fire;
  wire                when_CMemHost_l67;
  wire                io_hostd_bpss_rd_done_fire;
  wire                io_hostd_bpss_wr_done_fire;
  wire                when_CMemHost_l76;
  wire                io_hostd_axis_host_sink_fire;
  wire                io_hostd_axis_host_src_fire;
  wire                cmemToReq;
  wire                io_axi_cmem_aw_fire;
  wire                io_axi_cmem_ar_fire;
  wire                when_CMemHost_l116;
  wire                io_axi_cmem_aw_fire_1;
  wire                io_axi_cmem_ar_fire_1;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                when_CMemHost_l24;
  wire                when_CMemHost_l25;
  wire                when_CMemHost_l37;
  wire                when_CMemHost_l42;
  wire                when_StateMachine_l234;
  `ifndef SYNTHESIS
  reg [31:0] fsm_stateReg_string;
  reg [31:0] fsm_stateNext_string;
  `endif


  assign _zz_reqHostAddr = {48'd0, io_len};
  assign _zz_io_axi_cmem_aw_payload_len = (_zz_io_axi_cmem_aw_payload_len_1 - 10'h001);
  assign _zz_io_axi_cmem_aw_payload_len_1 = (io_len >>> 6);
  assign _zz_io_axi_cmem_ar_payload_len = (_zz_io_axi_cmem_ar_payload_len_1 - 10'h001);
  assign _zz_io_axi_cmem_ar_payload_len_1 = (io_len >>> 6);
  assign _zz_cmemWrAddr = {48'd0, io_len};
  assign _zz_cmemRdAddr = {48'd0, io_len};
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_BOOT : fsm_stateReg_string = "BOOT";
      fsm_enumDef_IDLE : fsm_stateReg_string = "IDLE";
      fsm_enumDef_RD : fsm_stateReg_string = "RD  ";
      fsm_enumDef_WR : fsm_stateReg_string = "WR  ";
      default : fsm_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_BOOT : fsm_stateNext_string = "BOOT";
      fsm_enumDef_IDLE : fsm_stateNext_string = "IDLE";
      fsm_enumDef_RD : fsm_stateNext_string = "RD  ";
      fsm_enumDef_WR : fsm_stateNext_string = "WR  ";
      default : fsm_stateNext_string = "????";
    endcase
  end
  `endif

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_RD : begin
      end
      fsm_enumDef_WR : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  assign bpss_rd_req_vaddr = reqHostAddr[47:0];
  assign bpss_rd_req_len = {12'd0, io_len};
  assign bpss_rd_req_stream = 1'b0;
  assign bpss_rd_req_sync = 1'b0;
  assign bpss_rd_req_ctl = 1'b1;
  assign bpss_rd_req_host = 1'b1;
  assign bpss_rd_req_dest = 4'b0000;
  assign bpss_rd_req_pid = io_pid;
  assign bpss_rd_req_vfid = 1'b0;
  assign bpss_rd_req_rsrvd = 5'h0;
  assign bpss_wr_req_vaddr = reqHostAddr[47:0];
  assign bpss_wr_req_len = {12'd0, io_len};
  assign bpss_wr_req_stream = 1'b0;
  assign bpss_wr_req_sync = 1'b0;
  assign bpss_wr_req_ctl = 1'b1;
  assign bpss_wr_req_host = 1'b1;
  assign bpss_wr_req_dest = 4'b0000;
  assign bpss_wr_req_pid = io_pid;
  assign bpss_wr_req_vfid = 1'b0;
  assign bpss_wr_req_rsrvd = 5'h0;
  assign io_hostd_bpss_rd_req_payload_data = {bpss_rd_req_vaddr,{bpss_rd_req_len,{bpss_rd_req_stream,{bpss_rd_req_sync,{bpss_rd_req_ctl,{bpss_rd_req_host,{bpss_rd_req_dest,{bpss_rd_req_pid,{bpss_rd_req_vfid,bpss_rd_req_rsrvd}}}}}}}}};
  assign io_hostd_bpss_wr_req_payload_data = {bpss_wr_req_vaddr,{bpss_wr_req_len,{bpss_wr_req_stream,{bpss_wr_req_sync,{bpss_wr_req_ctl,{bpss_wr_req_host,{bpss_wr_req_dest,{bpss_wr_req_pid,{bpss_wr_req_vfid,bpss_wr_req_rsrvd}}}}}}}}};
  assign io_hostd_bpss_rd_req_valid = ((cntHostReq != io_cnt) && (fsm_stateReg == fsm_enumDef_RD));
  assign io_hostd_bpss_wr_req_valid = ((cntHostReq != io_cnt) && (fsm_stateReg == fsm_enumDef_WR));
  assign io_hostd_bpss_rd_req_fire = (io_hostd_bpss_rd_req_valid && io_hostd_bpss_rd_req_ready);
  assign io_hostd_bpss_wr_req_fire = (io_hostd_bpss_wr_req_valid && io_hostd_bpss_wr_req_ready);
  assign when_CMemHost_l67 = (io_hostd_bpss_rd_req_fire || io_hostd_bpss_wr_req_fire);
  assign io_hostd_bpss_rd_done_ready = 1'b1;
  assign io_hostd_bpss_wr_done_ready = 1'b1;
  assign io_hostd_bpss_rd_done_fire = (io_hostd_bpss_rd_done_valid && io_hostd_bpss_rd_done_ready);
  assign io_hostd_bpss_wr_done_fire = (io_hostd_bpss_wr_done_valid && io_hostd_bpss_wr_done_ready);
  assign when_CMemHost_l76 = (io_hostd_bpss_rd_done_fire || io_hostd_bpss_wr_done_fire);
  assign io_hostd_axis_host_sink_fire = (io_hostd_axis_host_sink_valid && io_hostd_axis_host_sink_ready);
  assign io_hostd_axis_host_src_fire = (io_hostd_axis_host_src_valid && io_hostd_axis_host_src_ready);
  assign io_hostd_axis_host_src_payload_tdest = 4'b0000;
  assign io_hostd_axis_host_src_payload_tlast = 1'b0;
  assign io_hostd_axis_host_src_payload_tkeep = 64'hffffffffffffffff;
  assign io_axi_cmem_aw_payload_burst = 2'b01;
  assign io_axi_cmem_aw_payload_len = _zz_io_axi_cmem_aw_payload_len[7:0];
  assign io_axi_cmem_aw_payload_size = 3'b110;
  assign io_axi_cmem_aw_payload_addr = cmemWrAddr;
  assign io_axi_cmem_aw_payload_id = 6'h0;
  assign io_axi_cmem_w_payload_strb = 64'hffffffffffffffff;
  assign io_axi_cmem_w_payload_data = io_hostd_axis_host_sink_payload_tdata;
  assign io_axi_cmem_w_payload_last = io_hostd_axis_host_sink_payload_tlast;
  assign io_axi_cmem_w_valid = io_hostd_axis_host_sink_valid;
  assign io_hostd_axis_host_sink_ready = io_axi_cmem_w_ready;
  assign io_axi_cmem_b_ready = 1'b1;
  assign io_axi_cmem_ar_payload_burst = 2'b01;
  assign io_axi_cmem_ar_payload_len = _zz_io_axi_cmem_ar_payload_len[7:0];
  assign io_axi_cmem_ar_payload_size = 3'b110;
  assign io_axi_cmem_ar_payload_addr = cmemRdAddr;
  assign io_axi_cmem_ar_payload_id = 6'h0;
  assign io_hostd_axis_host_src_payload_tdata = io_axi_cmem_r_payload_data;
  assign io_hostd_axis_host_src_valid = io_axi_cmem_r_valid;
  assign io_axi_cmem_r_ready = io_hostd_axis_host_src_ready;
  assign cmemToReq = (cntHbmReq != io_cnt);
  assign io_axi_cmem_aw_valid = (cmemToReq && (fsm_stateReg == fsm_enumDef_RD));
  assign io_axi_cmem_ar_valid = (cmemToReq && (fsm_stateReg == fsm_enumDef_WR));
  assign io_axi_cmem_aw_fire = (io_axi_cmem_aw_valid && io_axi_cmem_aw_ready);
  assign io_axi_cmem_ar_fire = (io_axi_cmem_ar_valid && io_axi_cmem_ar_ready);
  assign when_CMemHost_l116 = (io_axi_cmem_aw_fire || io_axi_cmem_ar_fire);
  assign io_axi_cmem_aw_fire_1 = (io_axi_cmem_aw_valid && io_axi_cmem_aw_ready);
  assign io_axi_cmem_ar_fire_1 = (io_axi_cmem_ar_valid && io_axi_cmem_ar_ready);
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
        if(when_CMemHost_l24) begin
          fsm_stateNext = fsm_enumDef_RD;
        end
        if(when_CMemHost_l25) begin
          fsm_stateNext = fsm_enumDef_WR;
        end
      end
      fsm_enumDef_RD : begin
        if(when_CMemHost_l37) begin
          fsm_stateNext = fsm_enumDef_IDLE;
        end
      end
      fsm_enumDef_WR : begin
        if(when_CMemHost_l42) begin
          fsm_stateNext = fsm_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_IDLE;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_BOOT;
    end
  end

  assign when_CMemHost_l24 = (io_mode[0] ^ io_mode[1]);
  assign when_CMemHost_l25 = (io_mode[0] && io_mode[1]);
  assign when_CMemHost_l37 = (io_cntDone == io_cnt);
  assign when_CMemHost_l42 = (io_cntDone == io_cnt);
  assign when_StateMachine_l234 = ((fsm_stateReg == fsm_enumDef_IDLE) && (! (fsm_stateNext == fsm_enumDef_IDLE)));
  always @(posedge clk) begin
    if(!resetn) begin
      io_cntDone <= 64'h0;
      cntWrData <= 64'h0;
      cntRdData <= 64'h0;
      cntHostReq <= 64'h0;
      cntHbmReq <= 64'h0;
      cmemRdAddr <= 64'h0;
      cmemWrAddr <= 64'h0;
      reqHostAddr <= 64'h0;
      fsm_stateReg <= fsm_enumDef_BOOT;
    end else begin
      if(when_CMemHost_l67) begin
        cntHostReq <= (cntHostReq + 64'h0000000000000001);
        reqHostAddr <= (reqHostAddr + _zz_reqHostAddr);
      end
      if(when_CMemHost_l76) begin
        io_cntDone <= (io_cntDone + 64'h0000000000000001);
      end
      if(io_hostd_axis_host_sink_fire) begin
        cntRdData <= (cntRdData + 64'h0000000000000001);
      end
      if(io_hostd_axis_host_src_fire) begin
        cntWrData <= (cntWrData + 64'h0000000000000001);
      end
      if(when_CMemHost_l116) begin
        cntHbmReq <= (cntHbmReq + 64'h0000000000000001);
      end
      if(io_axi_cmem_aw_fire_1) begin
        cmemWrAddr <= (cmemWrAddr + _zz_cmemWrAddr);
      end
      if(io_axi_cmem_ar_fire_1) begin
        cmemRdAddr <= (cmemRdAddr + _zz_cmemRdAddr);
      end
      fsm_stateReg <= fsm_stateNext;
      if(when_StateMachine_l234) begin
        reqHostAddr <= io_hostAddr;
        cmemRdAddr <= io_cmemAddr;
        cmemWrAddr <= io_cmemAddr;
        cntRdData <= 64'h0;
        cntWrData <= 64'h0;
        cntHostReq <= 64'h0;
        cntHbmReq <= 64'h0;
        io_cntDone <= 64'h0;
      end
    end
  end


endmodule

module RdmaArb (
  output              io_rdmaV_0_rd_req_valid,
  input               io_rdmaV_0_rd_req_ready,
  output     [95:0]   io_rdmaV_0_rd_req_payload_data,
  output              io_rdmaV_0_wr_req_valid,
  input               io_rdmaV_0_wr_req_ready,
  output     [95:0]   io_rdmaV_0_wr_req_payload_data,
  input               io_rdmaV_0_sq_valid,
  output              io_rdmaV_0_sq_ready,
  input      [543:0]  io_rdmaV_0_sq_payload_data,
  output              io_rdmaV_0_ack_valid,
  input               io_rdmaV_0_ack_ready,
  output     [42:0]   io_rdmaV_0_ack_payload_data,
  output              io_rdmaV_0_axis_sink_valid,
  input               io_rdmaV_0_axis_sink_ready,
  output     [511:0]  io_rdmaV_0_axis_sink_payload_tdata,
  output     [63:0]   io_rdmaV_0_axis_sink_payload_tkeep,
  output              io_rdmaV_0_axis_sink_payload_tlast,
  input               io_rdmaV_0_axis_src_valid,
  output              io_rdmaV_0_axis_src_ready,
  input      [511:0]  io_rdmaV_0_axis_src_payload_tdata,
  input      [63:0]   io_rdmaV_0_axis_src_payload_tkeep,
  input               io_rdmaV_0_axis_src_payload_tlast,
  output              io_rdmaV_1_rd_req_valid,
  input               io_rdmaV_1_rd_req_ready,
  output     [95:0]   io_rdmaV_1_rd_req_payload_data,
  output              io_rdmaV_1_wr_req_valid,
  input               io_rdmaV_1_wr_req_ready,
  output     [95:0]   io_rdmaV_1_wr_req_payload_data,
  input               io_rdmaV_1_sq_valid,
  output              io_rdmaV_1_sq_ready,
  input      [543:0]  io_rdmaV_1_sq_payload_data,
  output              io_rdmaV_1_ack_valid,
  input               io_rdmaV_1_ack_ready,
  output     [42:0]   io_rdmaV_1_ack_payload_data,
  output              io_rdmaV_1_axis_sink_valid,
  input               io_rdmaV_1_axis_sink_ready,
  output     [511:0]  io_rdmaV_1_axis_sink_payload_tdata,
  output     [63:0]   io_rdmaV_1_axis_sink_payload_tkeep,
  output              io_rdmaV_1_axis_sink_payload_tlast,
  input               io_rdmaV_1_axis_src_valid,
  output              io_rdmaV_1_axis_src_ready,
  input      [511:0]  io_rdmaV_1_axis_src_payload_tdata,
  input      [63:0]   io_rdmaV_1_axis_src_payload_tkeep,
  input               io_rdmaV_1_axis_src_payload_tlast,
  input               io_rdmaio_rd_req_valid,
  output              io_rdmaio_rd_req_ready,
  input      [95:0]   io_rdmaio_rd_req_payload_data,
  input               io_rdmaio_wr_req_valid,
  output              io_rdmaio_wr_req_ready,
  input      [95:0]   io_rdmaio_wr_req_payload_data,
  output              io_rdmaio_sq_valid,
  input               io_rdmaio_sq_ready,
  output     [543:0]  io_rdmaio_sq_payload_data,
  input               io_rdmaio_ack_valid,
  output              io_rdmaio_ack_ready,
  input      [42:0]   io_rdmaio_ack_payload_data,
  input               io_rdmaio_axis_sink_valid,
  output              io_rdmaio_axis_sink_ready,
  input      [511:0]  io_rdmaio_axis_sink_payload_tdata,
  input      [63:0]   io_rdmaio_axis_sink_payload_tkeep,
  input               io_rdmaio_axis_sink_payload_tlast,
  output              io_rdmaio_axis_src_valid,
  input               io_rdmaio_axis_src_ready,
  output     [511:0]  io_rdmaio_axis_src_payload_tdata,
  output     [63:0]   io_rdmaio_axis_src_payload_tkeep,
  output              io_rdmaio_axis_src_payload_tlast,
  input               clk,
  input               resetn
);

  wire                strmFifo1_io_pop_ready;
  wire                strmFifo2_io_push_valid;
  wire                strmFifo2_io_pop_ready;
  wire                streamMux_2_io_output_ready;
  wire                streamDemux_7_io_input_valid;
  wire                streamMux_3_io_output_ready;
  wire                strmFifo3_io_pop_ready;
  wire                streamDemux_8_io_input_valid;
  wire                streamDemux_9_io_input_valid;
  wire       [0:0]    streamDemux_10_io_select;
  wire                strmFifo1_io_push_ready;
  wire                strmFifo1_io_pop_valid;
  wire       [0:0]    strmFifo1_io_pop_payload;
  wire       [5:0]    strmFifo1_io_occupancy;
  wire       [5:0]    strmFifo1_io_availability;
  wire                strmFifo2_io_push_ready;
  wire                strmFifo2_io_pop_valid;
  wire       [0:0]    strmFifo2_io_pop_payload;
  wire       [5:0]    strmFifo2_io_occupancy;
  wire       [5:0]    strmFifo2_io_availability;
  wire                streamMux_2_io_inputs_0_ready;
  wire                streamMux_2_io_inputs_1_ready;
  wire                streamMux_2_io_output_valid;
  wire       [543:0]  streamMux_2_io_output_payload_data;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [95:0]   streamDemux_7_io_outputs_0_payload_data;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [95:0]   streamDemux_7_io_outputs_1_payload_data;
  wire                streamMux_3_io_inputs_0_ready;
  wire                streamMux_3_io_inputs_1_ready;
  wire                streamMux_3_io_output_valid;
  wire       [511:0]  streamMux_3_io_output_payload_tdata;
  wire       [63:0]   streamMux_3_io_output_payload_tkeep;
  wire                streamMux_3_io_output_payload_tlast;
  wire                strmFifo3_io_push_ready;
  wire                strmFifo3_io_pop_valid;
  wire       [0:0]    strmFifo3_io_pop_payload;
  wire       [5:0]    strmFifo3_io_occupancy;
  wire       [5:0]    strmFifo3_io_availability;
  wire                streamDemux_8_io_input_ready;
  wire                streamDemux_8_io_outputs_0_valid;
  wire       [95:0]   streamDemux_8_io_outputs_0_payload_data;
  wire                streamDemux_8_io_outputs_1_valid;
  wire       [95:0]   streamDemux_8_io_outputs_1_payload_data;
  wire                streamDemux_9_io_input_ready;
  wire                streamDemux_9_io_outputs_0_valid;
  wire       [511:0]  streamDemux_9_io_outputs_0_payload_tdata;
  wire       [63:0]   streamDemux_9_io_outputs_0_payload_tkeep;
  wire                streamDemux_9_io_outputs_0_payload_tlast;
  wire                streamDemux_9_io_outputs_1_valid;
  wire       [511:0]  streamDemux_9_io_outputs_1_payload_tdata;
  wire       [63:0]   streamDemux_9_io_outputs_1_payload_tkeep;
  wire                streamDemux_9_io_outputs_1_payload_tlast;
  wire                streamDemux_10_io_input_ready;
  wire                streamDemux_10_io_outputs_0_valid;
  wire       [42:0]   streamDemux_10_io_outputs_0_payload_data;
  wire                streamDemux_10_io_outputs_1_valid;
  wire       [42:0]   streamDemux_10_io_outputs_1_payload_data;
  wire       [3:0]    _zz__zz_mskSqSel_2;
  wire       [3:0]    _zz__zz_mskSqSel_2_1;
  wire       [1:0]    _zz__zz_mskSqSel_2_2;
  wire       [9:0]    _zz_io_select;
  wire                sqV_0_valid;
  wire                sqV_0_ready;
  wire       [543:0]  sqV_0_payload_data;
  wire                sqV_1_valid;
  wire                sqV_1_ready;
  wire       [543:0]  sqV_1_payload_data;
  wire                io_rdmaV_0_sq_s2mPipe_valid;
  reg                 io_rdmaV_0_sq_s2mPipe_ready;
  wire       [543:0]  io_rdmaV_0_sq_s2mPipe_payload_data;
  reg                 io_rdmaV_0_sq_rValid;
  reg        [543:0]  io_rdmaV_0_sq_rData_data;
  wire                io_rdmaV_0_sq_s2mPipe_m2sPipe_valid;
  wire                io_rdmaV_0_sq_s2mPipe_m2sPipe_ready;
  wire       [543:0]  io_rdmaV_0_sq_s2mPipe_m2sPipe_payload_data;
  reg                 io_rdmaV_0_sq_s2mPipe_rValid;
  reg        [543:0]  io_rdmaV_0_sq_s2mPipe_rData_data;
  wire                when_Stream_l368;
  wire                io_rdmaV_1_sq_s2mPipe_valid;
  reg                 io_rdmaV_1_sq_s2mPipe_ready;
  wire       [543:0]  io_rdmaV_1_sq_s2mPipe_payload_data;
  reg                 io_rdmaV_1_sq_rValid;
  reg        [543:0]  io_rdmaV_1_sq_rData_data;
  wire                io_rdmaV_1_sq_s2mPipe_m2sPipe_valid;
  wire                io_rdmaV_1_sq_s2mPipe_m2sPipe_ready;
  wire       [543:0]  io_rdmaV_1_sq_s2mPipe_m2sPipe_payload_data;
  reg                 io_rdmaV_1_sq_s2mPipe_rValid;
  reg        [543:0]  io_rdmaV_1_sq_s2mPipe_rData_data;
  wire                when_Stream_l368_1;
  reg        [1:0]    mskSqVld;
  wire       [1:0]    mskSqSel;
  wire                io_rdmaio_sq_fire;
  reg        [1:0]    mskLocked;
  wire       [1:0]    _zz_mskSqSel;
  wire       [3:0]    _zz_mskSqSel_1;
  wire       [3:0]    _zz_mskSqSel_2;
  wire                _zz_sqSel;
  wire       [0:0]    sqSel;
  wire                _zz_io_rdmaio_sq_valid;
  wire                io_rdmaio_sq_fire_1;
  wire                io_rdmaio_rd_req_fire;
  wire                io_rdmaio_axis_src_fire;
  wire       [4:0]    wrReq_rsrvd;
  wire       [0:0]    wrReq_vfid;
  wire       [5:0]    wrReq_pid;
  wire       [3:0]    wrReq_dest;
  wire                wrReq_host;
  wire                wrReq_ctl;
  wire                wrReq_sync;
  wire                wrReq_stream;
  wire       [27:0]   wrReq_len;
  wire       [47:0]   wrReq_vaddr;
  wire       [0:0]    wrSel;
  wire                _zz_io_rdmaio_wr_req_ready;
  wire                io_rdmaio_wr_req_fire;
  wire                io_rdmaio_axis_sink_fire;

  assign _zz__zz_mskSqSel_2 = (_zz_mskSqSel_1 - _zz__zz_mskSqSel_2_1);
  assign _zz__zz_mskSqSel_2_2 = {mskLocked[0],mskLocked[1 : 1]};
  assign _zz__zz_mskSqSel_2_1 = {2'd0, _zz__zz_mskSqSel_2_2};
  assign _zz_io_select = io_rdmaio_ack_payload_data[10 : 1];
  StreamFifo_7 strmFifo1 (
    .io_push_valid   (io_rdmaio_sq_fire_1           ), //i
    .io_push_ready   (strmFifo1_io_push_ready       ), //o
    .io_push_payload (sqSel                         ), //i
    .io_pop_valid    (strmFifo1_io_pop_valid        ), //o
    .io_pop_ready    (strmFifo1_io_pop_ready        ), //i
    .io_pop_payload  (strmFifo1_io_pop_payload      ), //o
    .io_flush        (1'b0                          ), //i
    .io_occupancy    (strmFifo1_io_occupancy[5:0]   ), //o
    .io_availability (strmFifo1_io_availability[5:0]), //o
    .clk             (clk                           ), //i
    .resetn          (resetn                        )  //i
  );
  StreamFifo_7 strmFifo2 (
    .io_push_valid   (strmFifo2_io_push_valid       ), //i
    .io_push_ready   (strmFifo2_io_push_ready       ), //o
    .io_push_payload (strmFifo1_io_pop_payload      ), //i
    .io_pop_valid    (strmFifo2_io_pop_valid        ), //o
    .io_pop_ready    (strmFifo2_io_pop_ready        ), //i
    .io_pop_payload  (strmFifo2_io_pop_payload      ), //o
    .io_flush        (1'b0                          ), //i
    .io_occupancy    (strmFifo2_io_occupancy[5:0]   ), //o
    .io_availability (strmFifo2_io_availability[5:0]), //o
    .clk             (clk                           ), //i
    .resetn          (resetn                        )  //i
  );
  StreamMux streamMux_2 (
    .io_select                (sqSel                                    ), //i
    .io_inputs_0_valid        (sqV_0_valid                              ), //i
    .io_inputs_0_ready        (streamMux_2_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_data (sqV_0_payload_data[543:0]                ), //i
    .io_inputs_1_valid        (sqV_1_valid                              ), //i
    .io_inputs_1_ready        (streamMux_2_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_data (sqV_1_payload_data[543:0]                ), //i
    .io_output_valid          (streamMux_2_io_output_valid              ), //o
    .io_output_ready          (streamMux_2_io_output_ready              ), //i
    .io_output_payload_data   (streamMux_2_io_output_payload_data[543:0])  //o
  );
  StreamDemux_3 streamDemux_7 (
    .io_select                 (strmFifo1_io_pop_payload                     ), //i
    .io_input_valid            (streamDemux_7_io_input_valid                 ), //i
    .io_input_ready            (streamDemux_7_io_input_ready                 ), //o
    .io_input_payload_data     (io_rdmaio_rd_req_payload_data[95:0]          ), //i
    .io_outputs_0_valid        (streamDemux_7_io_outputs_0_valid             ), //o
    .io_outputs_0_ready        (io_rdmaV_0_rd_req_ready                      ), //i
    .io_outputs_0_payload_data (streamDemux_7_io_outputs_0_payload_data[95:0]), //o
    .io_outputs_1_valid        (streamDemux_7_io_outputs_1_valid             ), //o
    .io_outputs_1_ready        (io_rdmaV_1_rd_req_ready                      ), //i
    .io_outputs_1_payload_data (streamDemux_7_io_outputs_1_payload_data[95:0])  //o
  );
  StreamMux_1 streamMux_3 (
    .io_select                 (strmFifo2_io_pop_payload                  ), //i
    .io_inputs_0_valid         (io_rdmaV_0_axis_src_valid                 ), //i
    .io_inputs_0_ready         (streamMux_3_io_inputs_0_ready             ), //o
    .io_inputs_0_payload_tdata (io_rdmaV_0_axis_src_payload_tdata[511:0]  ), //i
    .io_inputs_0_payload_tkeep (io_rdmaV_0_axis_src_payload_tkeep[63:0]   ), //i
    .io_inputs_0_payload_tlast (io_rdmaV_0_axis_src_payload_tlast         ), //i
    .io_inputs_1_valid         (io_rdmaV_1_axis_src_valid                 ), //i
    .io_inputs_1_ready         (streamMux_3_io_inputs_1_ready             ), //o
    .io_inputs_1_payload_tdata (io_rdmaV_1_axis_src_payload_tdata[511:0]  ), //i
    .io_inputs_1_payload_tkeep (io_rdmaV_1_axis_src_payload_tkeep[63:0]   ), //i
    .io_inputs_1_payload_tlast (io_rdmaV_1_axis_src_payload_tlast         ), //i
    .io_output_valid           (streamMux_3_io_output_valid               ), //o
    .io_output_ready           (streamMux_3_io_output_ready               ), //i
    .io_output_payload_tdata   (streamMux_3_io_output_payload_tdata[511:0]), //o
    .io_output_payload_tkeep   (streamMux_3_io_output_payload_tkeep[63:0] ), //o
    .io_output_payload_tlast   (streamMux_3_io_output_payload_tlast       )  //o
  );
  StreamFifo_7 strmFifo3 (
    .io_push_valid   (io_rdmaio_wr_req_fire         ), //i
    .io_push_ready   (strmFifo3_io_push_ready       ), //o
    .io_push_payload (wrSel                         ), //i
    .io_pop_valid    (strmFifo3_io_pop_valid        ), //o
    .io_pop_ready    (strmFifo3_io_pop_ready        ), //i
    .io_pop_payload  (strmFifo3_io_pop_payload      ), //o
    .io_flush        (1'b0                          ), //i
    .io_occupancy    (strmFifo3_io_occupancy[5:0]   ), //o
    .io_availability (strmFifo3_io_availability[5:0]), //o
    .clk             (clk                           ), //i
    .resetn          (resetn                        )  //i
  );
  StreamDemux_3 streamDemux_8 (
    .io_select                 (wrSel                                        ), //i
    .io_input_valid            (streamDemux_8_io_input_valid                 ), //i
    .io_input_ready            (streamDemux_8_io_input_ready                 ), //o
    .io_input_payload_data     (io_rdmaio_wr_req_payload_data[95:0]          ), //i
    .io_outputs_0_valid        (streamDemux_8_io_outputs_0_valid             ), //o
    .io_outputs_0_ready        (io_rdmaV_0_wr_req_ready                      ), //i
    .io_outputs_0_payload_data (streamDemux_8_io_outputs_0_payload_data[95:0]), //o
    .io_outputs_1_valid        (streamDemux_8_io_outputs_1_valid             ), //o
    .io_outputs_1_ready        (io_rdmaV_1_wr_req_ready                      ), //i
    .io_outputs_1_payload_data (streamDemux_8_io_outputs_1_payload_data[95:0])  //o
  );
  StreamDemux_5 streamDemux_9 (
    .io_select                  (strmFifo3_io_pop_payload                       ), //i
    .io_input_valid             (streamDemux_9_io_input_valid                   ), //i
    .io_input_ready             (streamDemux_9_io_input_ready                   ), //o
    .io_input_payload_tdata     (io_rdmaio_axis_sink_payload_tdata[511:0]       ), //i
    .io_input_payload_tkeep     (io_rdmaio_axis_sink_payload_tkeep[63:0]        ), //i
    .io_input_payload_tlast     (io_rdmaio_axis_sink_payload_tlast              ), //i
    .io_outputs_0_valid         (streamDemux_9_io_outputs_0_valid               ), //o
    .io_outputs_0_ready         (io_rdmaV_0_axis_sink_ready                     ), //i
    .io_outputs_0_payload_tdata (streamDemux_9_io_outputs_0_payload_tdata[511:0]), //o
    .io_outputs_0_payload_tkeep (streamDemux_9_io_outputs_0_payload_tkeep[63:0] ), //o
    .io_outputs_0_payload_tlast (streamDemux_9_io_outputs_0_payload_tlast       ), //o
    .io_outputs_1_valid         (streamDemux_9_io_outputs_1_valid               ), //o
    .io_outputs_1_ready         (io_rdmaV_1_axis_sink_ready                     ), //i
    .io_outputs_1_payload_tdata (streamDemux_9_io_outputs_1_payload_tdata[511:0]), //o
    .io_outputs_1_payload_tkeep (streamDemux_9_io_outputs_1_payload_tkeep[63:0] ), //o
    .io_outputs_1_payload_tlast (streamDemux_9_io_outputs_1_payload_tlast       )  //o
  );
  StreamDemux_6 streamDemux_10 (
    .io_select                 (streamDemux_10_io_select                      ), //i
    .io_input_valid            (io_rdmaio_ack_valid                           ), //i
    .io_input_ready            (streamDemux_10_io_input_ready                 ), //o
    .io_input_payload_data     (io_rdmaio_ack_payload_data[42:0]              ), //i
    .io_outputs_0_valid        (streamDemux_10_io_outputs_0_valid             ), //o
    .io_outputs_0_ready        (io_rdmaV_0_ack_ready                          ), //i
    .io_outputs_0_payload_data (streamDemux_10_io_outputs_0_payload_data[42:0]), //o
    .io_outputs_1_valid        (streamDemux_10_io_outputs_1_valid             ), //o
    .io_outputs_1_ready        (io_rdmaV_1_ack_ready                          ), //i
    .io_outputs_1_payload_data (streamDemux_10_io_outputs_1_payload_data[42:0])  //o
  );
  assign io_rdmaV_0_sq_ready = (! io_rdmaV_0_sq_rValid);
  assign io_rdmaV_0_sq_s2mPipe_valid = (io_rdmaV_0_sq_valid || io_rdmaV_0_sq_rValid);
  assign io_rdmaV_0_sq_s2mPipe_payload_data = (io_rdmaV_0_sq_rValid ? io_rdmaV_0_sq_rData_data : io_rdmaV_0_sq_payload_data);
  always @(*) begin
    io_rdmaV_0_sq_s2mPipe_ready = io_rdmaV_0_sq_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      io_rdmaV_0_sq_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! io_rdmaV_0_sq_s2mPipe_m2sPipe_valid);
  assign io_rdmaV_0_sq_s2mPipe_m2sPipe_valid = io_rdmaV_0_sq_s2mPipe_rValid;
  assign io_rdmaV_0_sq_s2mPipe_m2sPipe_payload_data = io_rdmaV_0_sq_s2mPipe_rData_data;
  assign sqV_0_valid = io_rdmaV_0_sq_s2mPipe_m2sPipe_valid;
  assign io_rdmaV_0_sq_s2mPipe_m2sPipe_ready = sqV_0_ready;
  assign sqV_0_payload_data = io_rdmaV_0_sq_s2mPipe_m2sPipe_payload_data;
  assign io_rdmaV_1_sq_ready = (! io_rdmaV_1_sq_rValid);
  assign io_rdmaV_1_sq_s2mPipe_valid = (io_rdmaV_1_sq_valid || io_rdmaV_1_sq_rValid);
  assign io_rdmaV_1_sq_s2mPipe_payload_data = (io_rdmaV_1_sq_rValid ? io_rdmaV_1_sq_rData_data : io_rdmaV_1_sq_payload_data);
  always @(*) begin
    io_rdmaV_1_sq_s2mPipe_ready = io_rdmaV_1_sq_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      io_rdmaV_1_sq_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! io_rdmaV_1_sq_s2mPipe_m2sPipe_valid);
  assign io_rdmaV_1_sq_s2mPipe_m2sPipe_valid = io_rdmaV_1_sq_s2mPipe_rValid;
  assign io_rdmaV_1_sq_s2mPipe_m2sPipe_payload_data = io_rdmaV_1_sq_s2mPipe_rData_data;
  assign sqV_1_valid = io_rdmaV_1_sq_s2mPipe_m2sPipe_valid;
  assign io_rdmaV_1_sq_s2mPipe_m2sPipe_ready = sqV_1_ready;
  assign sqV_1_payload_data = io_rdmaV_1_sq_s2mPipe_m2sPipe_payload_data;
  always @(*) begin
    mskSqVld[0] = sqV_0_valid;
    mskSqVld[1] = sqV_1_valid;
  end

  assign io_rdmaio_sq_fire = (io_rdmaio_sq_valid && io_rdmaio_sq_ready);
  assign _zz_mskSqSel = mskSqVld;
  assign _zz_mskSqSel_1 = {_zz_mskSqSel,_zz_mskSqSel};
  assign _zz_mskSqSel_2 = (_zz_mskSqSel_1 & (~ _zz__zz_mskSqSel_2));
  assign mskSqSel = (_zz_mskSqSel_2[3 : 2] | _zz_mskSqSel_2[1 : 0]);
  assign _zz_sqSel = mskSqSel[1];
  assign sqSel = _zz_sqSel;
  assign sqV_0_ready = streamMux_2_io_inputs_0_ready;
  assign sqV_1_ready = streamMux_2_io_inputs_1_ready;
  assign _zz_io_rdmaio_sq_valid = (6'h0 < strmFifo1_io_availability);
  assign streamMux_2_io_output_ready = (io_rdmaio_sq_ready && _zz_io_rdmaio_sq_valid);
  assign io_rdmaio_sq_valid = (streamMux_2_io_output_valid && _zz_io_rdmaio_sq_valid);
  assign io_rdmaio_sq_payload_data = streamMux_2_io_output_payload_data;
  assign io_rdmaio_sq_fire_1 = (io_rdmaio_sq_valid && io_rdmaio_sq_ready);
  assign io_rdmaio_rd_req_ready = (streamDemux_7_io_input_ready && strmFifo1_io_pop_valid);
  assign streamDemux_7_io_input_valid = (io_rdmaio_rd_req_valid && strmFifo1_io_pop_valid);
  assign io_rdmaV_0_rd_req_valid = streamDemux_7_io_outputs_0_valid;
  assign io_rdmaV_0_rd_req_payload_data = streamDemux_7_io_outputs_0_payload_data;
  assign io_rdmaV_1_rd_req_valid = streamDemux_7_io_outputs_1_valid;
  assign io_rdmaV_1_rd_req_payload_data = streamDemux_7_io_outputs_1_payload_data;
  assign io_rdmaio_rd_req_fire = (io_rdmaio_rd_req_valid && io_rdmaio_rd_req_ready);
  assign strmFifo1_io_pop_ready = (strmFifo2_io_push_ready && io_rdmaio_rd_req_fire);
  assign strmFifo2_io_push_valid = (strmFifo1_io_pop_valid && io_rdmaio_rd_req_fire);
  assign io_rdmaV_0_axis_src_ready = streamMux_3_io_inputs_0_ready;
  assign io_rdmaV_1_axis_src_ready = streamMux_3_io_inputs_1_ready;
  assign streamMux_3_io_output_ready = (io_rdmaio_axis_src_ready && strmFifo2_io_pop_valid);
  assign io_rdmaio_axis_src_valid = (streamMux_3_io_output_valid && strmFifo2_io_pop_valid);
  assign io_rdmaio_axis_src_payload_tdata = streamMux_3_io_output_payload_tdata;
  assign io_rdmaio_axis_src_payload_tkeep = streamMux_3_io_output_payload_tkeep;
  assign io_rdmaio_axis_src_payload_tlast = streamMux_3_io_output_payload_tlast;
  assign io_rdmaio_axis_src_fire = (io_rdmaio_axis_src_valid && io_rdmaio_axis_src_ready);
  assign strmFifo2_io_pop_ready = (io_rdmaio_axis_src_fire && io_rdmaio_axis_src_payload_tlast);
  assign wrReq_rsrvd = io_rdmaio_wr_req_payload_data[4 : 0];
  assign wrReq_vfid = io_rdmaio_wr_req_payload_data[5 : 5];
  assign wrReq_pid = io_rdmaio_wr_req_payload_data[11 : 6];
  assign wrReq_dest = io_rdmaio_wr_req_payload_data[15 : 12];
  assign wrReq_host = io_rdmaio_wr_req_payload_data[16];
  assign wrReq_ctl = io_rdmaio_wr_req_payload_data[17];
  assign wrReq_sync = io_rdmaio_wr_req_payload_data[18];
  assign wrReq_stream = io_rdmaio_wr_req_payload_data[19];
  assign wrReq_len = io_rdmaio_wr_req_payload_data[47 : 20];
  assign wrReq_vaddr = io_rdmaio_wr_req_payload_data[95 : 48];
  assign wrSel = wrReq_vaddr[0:0];
  assign _zz_io_rdmaio_wr_req_ready = (6'h0 < strmFifo3_io_availability);
  assign io_rdmaio_wr_req_ready = (streamDemux_8_io_input_ready && _zz_io_rdmaio_wr_req_ready);
  assign streamDemux_8_io_input_valid = (io_rdmaio_wr_req_valid && _zz_io_rdmaio_wr_req_ready);
  assign io_rdmaV_0_wr_req_valid = streamDemux_8_io_outputs_0_valid;
  assign io_rdmaV_0_wr_req_payload_data = streamDemux_8_io_outputs_0_payload_data;
  assign io_rdmaV_1_wr_req_valid = streamDemux_8_io_outputs_1_valid;
  assign io_rdmaV_1_wr_req_payload_data = streamDemux_8_io_outputs_1_payload_data;
  assign io_rdmaio_wr_req_fire = (io_rdmaio_wr_req_valid && io_rdmaio_wr_req_ready);
  assign io_rdmaio_axis_sink_ready = (streamDemux_9_io_input_ready && strmFifo3_io_pop_valid);
  assign streamDemux_9_io_input_valid = (io_rdmaio_axis_sink_valid && strmFifo3_io_pop_valid);
  assign io_rdmaV_0_axis_sink_valid = streamDemux_9_io_outputs_0_valid;
  assign io_rdmaV_0_axis_sink_payload_tdata = streamDemux_9_io_outputs_0_payload_tdata;
  assign io_rdmaV_0_axis_sink_payload_tkeep = streamDemux_9_io_outputs_0_payload_tkeep;
  assign io_rdmaV_0_axis_sink_payload_tlast = streamDemux_9_io_outputs_0_payload_tlast;
  assign io_rdmaV_1_axis_sink_valid = streamDemux_9_io_outputs_1_valid;
  assign io_rdmaV_1_axis_sink_payload_tdata = streamDemux_9_io_outputs_1_payload_tdata;
  assign io_rdmaV_1_axis_sink_payload_tkeep = streamDemux_9_io_outputs_1_payload_tkeep;
  assign io_rdmaV_1_axis_sink_payload_tlast = streamDemux_9_io_outputs_1_payload_tlast;
  assign io_rdmaio_axis_sink_fire = (io_rdmaio_axis_sink_valid && io_rdmaio_axis_sink_ready);
  assign strmFifo3_io_pop_ready = (io_rdmaio_axis_sink_fire && io_rdmaio_axis_sink_payload_tlast);
  assign io_rdmaio_ack_ready = streamDemux_10_io_input_ready;
  assign streamDemux_10_io_select = _zz_io_select[0:0];
  assign io_rdmaV_0_ack_valid = streamDemux_10_io_outputs_0_valid;
  assign io_rdmaV_0_ack_payload_data = streamDemux_10_io_outputs_0_payload_data;
  assign io_rdmaV_1_ack_valid = streamDemux_10_io_outputs_1_valid;
  assign io_rdmaV_1_ack_payload_data = streamDemux_10_io_outputs_1_payload_data;
  always @(posedge clk) begin
    if(!resetn) begin
      io_rdmaV_0_sq_rValid <= 1'b0;
      io_rdmaV_0_sq_s2mPipe_rValid <= 1'b0;
      io_rdmaV_1_sq_rValid <= 1'b0;
      io_rdmaV_1_sq_s2mPipe_rValid <= 1'b0;
      mskLocked <= 2'b01;
    end else begin
      if(io_rdmaV_0_sq_valid) begin
        io_rdmaV_0_sq_rValid <= 1'b1;
      end
      if(io_rdmaV_0_sq_s2mPipe_ready) begin
        io_rdmaV_0_sq_rValid <= 1'b0;
      end
      if(io_rdmaV_0_sq_s2mPipe_ready) begin
        io_rdmaV_0_sq_s2mPipe_rValid <= io_rdmaV_0_sq_s2mPipe_valid;
      end
      if(io_rdmaV_1_sq_valid) begin
        io_rdmaV_1_sq_rValid <= 1'b1;
      end
      if(io_rdmaV_1_sq_s2mPipe_ready) begin
        io_rdmaV_1_sq_rValid <= 1'b0;
      end
      if(io_rdmaV_1_sq_s2mPipe_ready) begin
        io_rdmaV_1_sq_s2mPipe_rValid <= io_rdmaV_1_sq_s2mPipe_valid;
      end
      if(io_rdmaio_sq_fire) begin
        mskLocked <= mskSqSel;
      end
    end
  end

  always @(posedge clk) begin
    if(io_rdmaV_0_sq_ready) begin
      io_rdmaV_0_sq_rData_data <= io_rdmaV_0_sq_payload_data;
    end
    if(io_rdmaV_0_sq_s2mPipe_ready) begin
      io_rdmaV_0_sq_s2mPipe_rData_data <= io_rdmaV_0_sq_s2mPipe_payload_data;
    end
    if(io_rdmaV_1_sq_ready) begin
      io_rdmaV_1_sq_rData_data <= io_rdmaV_1_sq_payload_data;
    end
    if(io_rdmaV_1_sq_s2mPipe_ready) begin
      io_rdmaV_1_sq_s2mPipe_rData_data <= io_rdmaV_1_sq_s2mPipe_payload_data;
    end
  end


endmodule

module RdmaFlowBpss_1 (
  input               io_rdma_rd_req_valid,
  output              io_rdma_rd_req_ready,
  input      [95:0]   io_rdma_rd_req_payload_data,
  input               io_rdma_wr_req_valid,
  output              io_rdma_wr_req_ready,
  input      [95:0]   io_rdma_wr_req_payload_data,
  output              io_rdma_sq_valid,
  input               io_rdma_sq_ready,
  output     [543:0]  io_rdma_sq_payload_data,
  input               io_rdma_ack_valid,
  output              io_rdma_ack_ready,
  input      [42:0]   io_rdma_ack_payload_data,
  input               io_rdma_axis_sink_valid,
  output              io_rdma_axis_sink_ready,
  input      [511:0]  io_rdma_axis_sink_payload_tdata,
  input      [63:0]   io_rdma_axis_sink_payload_tkeep,
  input               io_rdma_axis_sink_payload_tlast,
  output              io_rdma_axis_src_valid,
  input               io_rdma_axis_src_ready,
  output     [511:0]  io_rdma_axis_src_payload_tdata,
  output     [63:0]   io_rdma_axis_src_payload_tkeep,
  output reg          io_rdma_axis_src_payload_tlast,
  input               io_q_sink_valid,
  output              io_q_sink_ready,
  input      [511:0]  io_q_sink_payload,
  output              io_q_src_valid,
  input               io_q_src_ready,
  output     [511:0]  io_q_src_payload,
  input               io_ctrl_en,
  input      [31:0]   io_ctrl_len,
  input      [9:0]    io_ctrl_qpn,
  input      [3:0]    io_ctrl_flowId,
  input               clk,
  input               resetn
);

  wire                streamFifo_10_io_flush;
  wire                streamFifo_11_io_pop_ready;
  wire                streamFifo_11_io_flush;
  wire                streamFifo_10_io_push_ready;
  wire                streamFifo_10_io_pop_valid;
  wire       [511:0]  streamFifo_10_io_pop_payload;
  wire       [9:0]    streamFifo_10_io_occupancy;
  wire       [9:0]    streamFifo_10_io_availability;
  wire                streamFifo_11_io_push_ready;
  wire                streamFifo_11_io_pop_valid;
  wire       [511:0]  streamFifo_11_io_pop_payload;
  wire       [9:0]    streamFifo_11_io_occupancy;
  wire       [9:0]    streamFifo_11_io_availability;
  wire       [8:0]    _zz__zz_io_rdma_sq_valid_2;
  wire       [0:0]    _zz__zz_io_rdma_sq_valid_2_1;
  wire       [25:0]   _zz_when_RdmaFlowBpss_l47_1;
  wire       [25:0]   _zz_when_RdmaFlowBpss_l47_2;
  wire       [11:0]   _zz_io_rdma_sq_valid_5;
  wire       [11:0]   _zz_io_rdma_sq_valid_6;
  wire       [11:0]   _zz_io_rdma_sq_valid_7;
  wire       [11:0]   _zz_io_rdma_sq_valid_8;
  wire       [11:0]   _zz_io_rdma_sq_valid_9;
  wire                incCntToSend;
  wire                io_rdma_axis_src_fire;
  wire                decCntToSend;
  reg        [7:0]    _zz_io_rdma_sq_valid;
  reg                 when_Utils_l21;
  wire       [1:0]    switch_Utils_l16;
  wire                timeOutInc;
  wire                io_rdma_sq_fire;
  wire                when_Utils_l63;
  reg                 _zz_io_rdma_sq_valid_1;
  reg                 _zz_1;
  reg        [8:0]    _zz_io_rdma_sq_valid_2;
  reg        [8:0]    _zz_io_rdma_sq_valid_3;
  wire                _zz_io_rdma_sq_valid_4;
  reg                 _zz_when_Utils_l65;
  wire                when_Utils_l65;
  wire                io_rdma_sq_fire_1;
  wire                when_RdmaFlowBpss_l44;
  reg                 rTimeOut;
  wire                io_rdma_axis_src_fire_1;
  reg        [25:0]   _zz_when_RdmaFlowBpss_l47;
  wire                when_RdmaFlowBpss_l47;
  reg                 _zz_when_Utils_l39;
  wire       [1:0]    switch_Utils_l34;
  wire                when_Utils_l39;
  wire       [63:0]   rdma_base_lvaddr;
  wire       [63:0]   rdma_base_rvaddr;
  wire       [31:0]   rdma_base_len;
  wire       [351:0]  rdma_base_params;
  wire       [13:0]   sq_rsrvd;
  wire       [511:0]  sq_msg;
  wire                sq_last;
  wire                sq_mode;
  wire                sq_host;
  wire       [9:0]    sq_qpn;
  wire       [4:0]    sq_opcode;
  wire                _zz_io_rdma_axis_src_valid;
  wire                when_RdmaFlowBpss_l117;

  assign _zz__zz_io_rdma_sq_valid_2_1 = _zz_io_rdma_sq_valid_1;
  assign _zz__zz_io_rdma_sq_valid_2 = {8'd0, _zz__zz_io_rdma_sq_valid_2_1};
  assign _zz_when_RdmaFlowBpss_l47_1 = ((rTimeOut ? 26'h0000001 : _zz_when_RdmaFlowBpss_l47_2) - 26'h0000001);
  assign _zz_when_RdmaFlowBpss_l47_2 = (io_ctrl_len >>> 6);
  assign _zz_io_rdma_sq_valid_5 = 12'h010;
  assign _zz_io_rdma_sq_valid_6 = _zz_io_rdma_sq_valid_7;
  assign _zz_io_rdma_sq_valid_7 = (_zz_io_rdma_sq_valid_8 - _zz_io_rdma_sq_valid_9);
  assign _zz_io_rdma_sq_valid_8 = {2'd0, streamFifo_11_io_occupancy};
  assign _zz_io_rdma_sq_valid_9 = ({4'd0,_zz_io_rdma_sq_valid} <<< 4);
  StreamFifo_3 streamFifo_10 (
    .io_push_valid   (io_rdma_axis_sink_valid               ), //i
    .io_push_ready   (streamFifo_10_io_push_ready           ), //o
    .io_push_payload (io_rdma_axis_sink_payload_tdata[511:0]), //i
    .io_pop_valid    (streamFifo_10_io_pop_valid            ), //o
    .io_pop_ready    (io_q_src_ready                        ), //i
    .io_pop_payload  (streamFifo_10_io_pop_payload[511:0]   ), //o
    .io_flush        (streamFifo_10_io_flush                ), //i
    .io_occupancy    (streamFifo_10_io_occupancy[9:0]       ), //o
    .io_availability (streamFifo_10_io_availability[9:0]    ), //o
    .clk             (clk                                   ), //i
    .resetn          (resetn                                )  //i
  );
  StreamFifo_3 streamFifo_11 (
    .io_push_valid   (io_q_sink_valid                    ), //i
    .io_push_ready   (streamFifo_11_io_push_ready        ), //o
    .io_push_payload (io_q_sink_payload[511:0]           ), //i
    .io_pop_valid    (streamFifo_11_io_pop_valid         ), //o
    .io_pop_ready    (streamFifo_11_io_pop_ready         ), //i
    .io_pop_payload  (streamFifo_11_io_pop_payload[511:0]), //o
    .io_flush        (streamFifo_11_io_flush             ), //i
    .io_occupancy    (streamFifo_11_io_occupancy[9:0]    ), //o
    .io_availability (streamFifo_11_io_availability[9:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  always @(*) begin
    io_rdma_axis_src_payload_tlast = 1'b0;
    if(when_RdmaFlowBpss_l47) begin
      io_rdma_axis_src_payload_tlast = 1'b1;
    end
  end

  assign io_rdma_axis_src_payload_tkeep = 64'hffffffffffffffff;
  assign io_rdma_ack_ready = 1'b1;
  assign io_rdma_rd_req_ready = 1'b1;
  assign io_rdma_wr_req_ready = 1'b1;
  assign incCntToSend = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign io_rdma_axis_src_fire = (io_rdma_axis_src_valid && io_rdma_axis_src_ready);
  assign decCntToSend = (io_rdma_axis_src_fire && io_rdma_axis_src_payload_tlast);
  always @(*) begin
    when_Utils_l21 = 1'b0;
    if(when_RdmaFlowBpss_l117) begin
      when_Utils_l21 = 1'b1;
    end
  end

  assign switch_Utils_l16 = {incCntToSend,decCntToSend};
  assign io_rdma_sq_fire = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign when_Utils_l63 = 1'b0;
  always @(*) begin
    _zz_io_rdma_sq_valid_1 = 1'b0;
    if(when_Utils_l65) begin
      _zz_io_rdma_sq_valid_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(io_rdma_sq_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_io_rdma_sq_valid_4 = (_zz_io_rdma_sq_valid_3 == 9'h1ff);
  always @(*) begin
    _zz_io_rdma_sq_valid_2 = (_zz_io_rdma_sq_valid_3 + _zz__zz_io_rdma_sq_valid_2);
    if(_zz_1) begin
      _zz_io_rdma_sq_valid_2 = 9'h0;
    end
  end

  assign when_Utils_l65 = ((timeOutInc && (! _zz_when_Utils_l65)) && (! _zz_io_rdma_sq_valid_4));
  assign io_rdma_sq_fire_1 = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign when_RdmaFlowBpss_l44 = (io_rdma_sq_fire_1 || decCntToSend);
  assign io_rdma_axis_src_fire_1 = (io_rdma_axis_src_valid && io_rdma_axis_src_ready);
  assign when_RdmaFlowBpss_l47 = (_zz_when_RdmaFlowBpss_l47 == _zz_when_RdmaFlowBpss_l47_1);
  always @(*) begin
    _zz_when_Utils_l39 = 1'b0;
    if(when_RdmaFlowBpss_l117) begin
      _zz_when_Utils_l39 = 1'b1;
    end
  end

  assign switch_Utils_l34 = {io_rdma_axis_src_fire_1,1'b0};
  assign when_Utils_l39 = (_zz_when_Utils_l39 || (when_RdmaFlowBpss_l47 && io_rdma_axis_src_fire_1));
  assign rdma_base_lvaddr = 64'h0;
  assign rdma_base_rvaddr = {60'd0, io_ctrl_flowId};
  assign rdma_base_len = (rTimeOut ? 32'h00000040 : io_ctrl_len);
  assign rdma_base_params = 352'h0;
  assign sq_opcode = 5'h0a;
  assign sq_qpn = io_ctrl_qpn;
  assign sq_host = 1'b0;
  assign sq_mode = 1'b1;
  assign sq_last = 1'b1;
  assign sq_msg = {rdma_base_params,{rdma_base_len,{rdma_base_rvaddr,rdma_base_lvaddr}}};
  assign sq_rsrvd = 14'h0;
  assign io_rdma_sq_payload_data = {sq_opcode,{sq_qpn,{sq_host,{sq_mode,{sq_last,{sq_msg,sq_rsrvd}}}}}};
  assign streamFifo_10_io_flush = (! io_ctrl_en);
  assign streamFifo_11_io_flush = (! io_ctrl_en);
  assign io_q_src_valid = streamFifo_10_io_pop_valid;
  assign io_q_src_payload = streamFifo_10_io_pop_payload;
  assign io_rdma_axis_sink_ready = streamFifo_10_io_push_ready;
  assign io_q_sink_ready = streamFifo_11_io_push_ready;
  assign _zz_io_rdma_axis_src_valid = (8'h0 < _zz_io_rdma_sq_valid);
  assign streamFifo_11_io_pop_ready = (io_rdma_axis_src_ready && _zz_io_rdma_axis_src_valid);
  assign io_rdma_axis_src_valid = (streamFifo_11_io_pop_valid && _zz_io_rdma_axis_src_valid);
  assign io_rdma_axis_src_payload_tdata = streamFifo_11_io_pop_payload;
  assign timeOutInc = (10'h0 < streamFifo_11_io_occupancy);
  assign io_rdma_sq_valid = (($signed(_zz_io_rdma_sq_valid_5) <= $signed(_zz_io_rdma_sq_valid_6)) || _zz_io_rdma_sq_valid_4);
  assign when_RdmaFlowBpss_l117 = (! io_ctrl_en);
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_rdma_sq_valid <= 8'h0;
      _zz_io_rdma_sq_valid_3 <= 9'h0;
      _zz_when_RdmaFlowBpss_l47 <= 26'h0;
    end else begin
      if((switch_Utils_l16 == {1'b1,1'b0})) begin
          _zz_io_rdma_sq_valid <= (_zz_io_rdma_sq_valid + 8'h01);
      end else if((switch_Utils_l16 == {1'b0,1'b1})) begin
          _zz_io_rdma_sq_valid <= (_zz_io_rdma_sq_valid - 8'h01);
      end
      if(when_Utils_l21) begin
        _zz_io_rdma_sq_valid <= 8'h0;
      end
      _zz_io_rdma_sq_valid_3 <= _zz_io_rdma_sq_valid_2;
      if((switch_Utils_l34 == {1'b1,1'b0})) begin
          _zz_when_RdmaFlowBpss_l47 <= (_zz_when_RdmaFlowBpss_l47 + 26'h0000001);
      end else if((switch_Utils_l34 == {1'b0,1'b1})) begin
          _zz_when_RdmaFlowBpss_l47 <= (_zz_when_RdmaFlowBpss_l47 - 26'h0000001);
      end
      if(when_Utils_l39) begin
        _zz_when_RdmaFlowBpss_l47 <= 26'h0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_Utils_l63) begin
      _zz_when_Utils_l65 <= 1'b1;
    end
    if(io_rdma_sq_fire) begin
      _zz_when_Utils_l65 <= 1'b0;
    end
    if(when_RdmaFlowBpss_l44) begin
      rTimeOut <= _zz_io_rdma_sq_valid_4;
    end
  end


endmodule

module RdmaFlowBpss (
  input               io_rdma_rd_req_valid,
  output              io_rdma_rd_req_ready,
  input      [95:0]   io_rdma_rd_req_payload_data,
  input               io_rdma_wr_req_valid,
  output              io_rdma_wr_req_ready,
  input      [95:0]   io_rdma_wr_req_payload_data,
  output              io_rdma_sq_valid,
  input               io_rdma_sq_ready,
  output     [543:0]  io_rdma_sq_payload_data,
  input               io_rdma_ack_valid,
  output              io_rdma_ack_ready,
  input      [42:0]   io_rdma_ack_payload_data,
  input               io_rdma_axis_sink_valid,
  output              io_rdma_axis_sink_ready,
  input      [511:0]  io_rdma_axis_sink_payload_tdata,
  input      [63:0]   io_rdma_axis_sink_payload_tkeep,
  input               io_rdma_axis_sink_payload_tlast,
  output              io_rdma_axis_src_valid,
  input               io_rdma_axis_src_ready,
  output     [511:0]  io_rdma_axis_src_payload_tdata,
  output     [63:0]   io_rdma_axis_src_payload_tkeep,
  output reg          io_rdma_axis_src_payload_tlast,
  input               io_q_sink_valid,
  output              io_q_sink_ready,
  input      [511:0]  io_q_sink_payload,
  output              io_q_src_valid,
  input               io_q_src_ready,
  output     [511:0]  io_q_src_payload,
  input               io_ctrl_en,
  input      [31:0]   io_ctrl_len,
  input      [9:0]    io_ctrl_qpn,
  input      [3:0]    io_ctrl_flowId,
  input               clk,
  input               resetn
);

  wire                streamFifo_10_io_pop_ready;
  wire                streamFifo_10_io_flush;
  wire                streamFifo_11_io_flush;
  wire                streamFifo_10_io_push_ready;
  wire                streamFifo_10_io_pop_valid;
  wire       [511:0]  streamFifo_10_io_pop_payload;
  wire       [9:0]    streamFifo_10_io_occupancy;
  wire       [9:0]    streamFifo_10_io_availability;
  wire                streamFifo_11_io_push_ready;
  wire                streamFifo_11_io_pop_valid;
  wire       [511:0]  streamFifo_11_io_pop_payload;
  wire       [9:0]    streamFifo_11_io_occupancy;
  wire       [9:0]    streamFifo_11_io_availability;
  wire       [8:0]    _zz__zz_io_rdma_sq_valid_2;
  wire       [0:0]    _zz__zz_io_rdma_sq_valid_2_1;
  wire       [25:0]   _zz_when_RdmaFlowBpss_l47_1;
  wire       [25:0]   _zz_when_RdmaFlowBpss_l47_2;
  wire       [11:0]   _zz_io_rdma_sq_valid_5;
  wire       [11:0]   _zz_io_rdma_sq_valid_6;
  wire       [11:0]   _zz_io_rdma_sq_valid_7;
  wire       [11:0]   _zz_io_rdma_sq_valid_8;
  wire       [11:0]   _zz_io_rdma_sq_valid_9;
  wire                incCntToSend;
  wire                io_rdma_axis_src_fire;
  wire                decCntToSend;
  reg        [7:0]    _zz_io_rdma_sq_valid;
  reg                 when_Utils_l21;
  wire       [1:0]    switch_Utils_l16;
  wire                timeOutInc;
  wire                io_rdma_sq_fire;
  wire                when_Utils_l63;
  reg                 _zz_io_rdma_sq_valid_1;
  reg                 _zz_1;
  reg        [8:0]    _zz_io_rdma_sq_valid_2;
  reg        [8:0]    _zz_io_rdma_sq_valid_3;
  wire                _zz_io_rdma_sq_valid_4;
  reg                 _zz_when_Utils_l65;
  wire                when_Utils_l65;
  wire                io_rdma_sq_fire_1;
  wire                when_RdmaFlowBpss_l44;
  reg                 rTimeOut;
  wire                io_rdma_axis_src_fire_1;
  reg        [25:0]   _zz_when_RdmaFlowBpss_l47;
  wire                when_RdmaFlowBpss_l47;
  reg                 _zz_when_Utils_l39;
  wire       [1:0]    switch_Utils_l34;
  wire                when_Utils_l39;
  wire       [63:0]   rdma_base_lvaddr;
  wire       [63:0]   rdma_base_rvaddr;
  wire       [31:0]   rdma_base_len;
  wire       [351:0]  rdma_base_params;
  wire       [13:0]   sq_rsrvd;
  wire       [511:0]  sq_msg;
  wire                sq_last;
  wire                sq_mode;
  wire                sq_host;
  wire       [9:0]    sq_qpn;
  wire       [4:0]    sq_opcode;
  wire                _zz_io_rdma_axis_src_valid;
  wire                when_RdmaFlowBpss_l117;

  assign _zz__zz_io_rdma_sq_valid_2_1 = _zz_io_rdma_sq_valid_1;
  assign _zz__zz_io_rdma_sq_valid_2 = {8'd0, _zz__zz_io_rdma_sq_valid_2_1};
  assign _zz_when_RdmaFlowBpss_l47_1 = ((rTimeOut ? 26'h0000001 : _zz_when_RdmaFlowBpss_l47_2) - 26'h0000001);
  assign _zz_when_RdmaFlowBpss_l47_2 = (io_ctrl_len >>> 6);
  assign _zz_io_rdma_sq_valid_5 = 12'h010;
  assign _zz_io_rdma_sq_valid_6 = _zz_io_rdma_sq_valid_7;
  assign _zz_io_rdma_sq_valid_7 = (_zz_io_rdma_sq_valid_8 - _zz_io_rdma_sq_valid_9);
  assign _zz_io_rdma_sq_valid_8 = {2'd0, streamFifo_10_io_occupancy};
  assign _zz_io_rdma_sq_valid_9 = ({4'd0,_zz_io_rdma_sq_valid} <<< 4);
  StreamFifo_3 streamFifo_10 (
    .io_push_valid   (io_q_sink_valid                    ), //i
    .io_push_ready   (streamFifo_10_io_push_ready        ), //o
    .io_push_payload (io_q_sink_payload[511:0]           ), //i
    .io_pop_valid    (streamFifo_10_io_pop_valid         ), //o
    .io_pop_ready    (streamFifo_10_io_pop_ready         ), //i
    .io_pop_payload  (streamFifo_10_io_pop_payload[511:0]), //o
    .io_flush        (streamFifo_10_io_flush             ), //i
    .io_occupancy    (streamFifo_10_io_occupancy[9:0]    ), //o
    .io_availability (streamFifo_10_io_availability[9:0] ), //o
    .clk             (clk                                ), //i
    .resetn          (resetn                             )  //i
  );
  StreamFifo_3 streamFifo_11 (
    .io_push_valid   (io_rdma_axis_sink_valid               ), //i
    .io_push_ready   (streamFifo_11_io_push_ready           ), //o
    .io_push_payload (io_rdma_axis_sink_payload_tdata[511:0]), //i
    .io_pop_valid    (streamFifo_11_io_pop_valid            ), //o
    .io_pop_ready    (io_q_src_ready                        ), //i
    .io_pop_payload  (streamFifo_11_io_pop_payload[511:0]   ), //o
    .io_flush        (streamFifo_11_io_flush                ), //i
    .io_occupancy    (streamFifo_11_io_occupancy[9:0]       ), //o
    .io_availability (streamFifo_11_io_availability[9:0]    ), //o
    .clk             (clk                                   ), //i
    .resetn          (resetn                                )  //i
  );
  always @(*) begin
    io_rdma_axis_src_payload_tlast = 1'b0;
    if(when_RdmaFlowBpss_l47) begin
      io_rdma_axis_src_payload_tlast = 1'b1;
    end
  end

  assign io_rdma_axis_src_payload_tkeep = 64'hffffffffffffffff;
  assign io_rdma_ack_ready = 1'b1;
  assign io_rdma_rd_req_ready = 1'b1;
  assign io_rdma_wr_req_ready = 1'b1;
  assign incCntToSend = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign io_rdma_axis_src_fire = (io_rdma_axis_src_valid && io_rdma_axis_src_ready);
  assign decCntToSend = (io_rdma_axis_src_fire && io_rdma_axis_src_payload_tlast);
  always @(*) begin
    when_Utils_l21 = 1'b0;
    if(when_RdmaFlowBpss_l117) begin
      when_Utils_l21 = 1'b1;
    end
  end

  assign switch_Utils_l16 = {incCntToSend,decCntToSend};
  assign io_rdma_sq_fire = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign when_Utils_l63 = 1'b0;
  always @(*) begin
    _zz_io_rdma_sq_valid_1 = 1'b0;
    if(when_Utils_l65) begin
      _zz_io_rdma_sq_valid_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(io_rdma_sq_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign _zz_io_rdma_sq_valid_4 = (_zz_io_rdma_sq_valid_3 == 9'h1ff);
  always @(*) begin
    _zz_io_rdma_sq_valid_2 = (_zz_io_rdma_sq_valid_3 + _zz__zz_io_rdma_sq_valid_2);
    if(_zz_1) begin
      _zz_io_rdma_sq_valid_2 = 9'h0;
    end
  end

  assign when_Utils_l65 = ((timeOutInc && (! _zz_when_Utils_l65)) && (! _zz_io_rdma_sq_valid_4));
  assign io_rdma_sq_fire_1 = (io_rdma_sq_valid && io_rdma_sq_ready);
  assign when_RdmaFlowBpss_l44 = (io_rdma_sq_fire_1 || decCntToSend);
  assign io_rdma_axis_src_fire_1 = (io_rdma_axis_src_valid && io_rdma_axis_src_ready);
  assign when_RdmaFlowBpss_l47 = (_zz_when_RdmaFlowBpss_l47 == _zz_when_RdmaFlowBpss_l47_1);
  always @(*) begin
    _zz_when_Utils_l39 = 1'b0;
    if(when_RdmaFlowBpss_l117) begin
      _zz_when_Utils_l39 = 1'b1;
    end
  end

  assign switch_Utils_l34 = {io_rdma_axis_src_fire_1,1'b0};
  assign when_Utils_l39 = (_zz_when_Utils_l39 || (when_RdmaFlowBpss_l47 && io_rdma_axis_src_fire_1));
  assign rdma_base_lvaddr = 64'h0;
  assign rdma_base_rvaddr = {60'd0, io_ctrl_flowId};
  assign rdma_base_len = (rTimeOut ? 32'h00000040 : io_ctrl_len);
  assign rdma_base_params = 352'h0;
  assign sq_opcode = 5'h0a;
  assign sq_qpn = io_ctrl_qpn;
  assign sq_host = 1'b0;
  assign sq_mode = 1'b1;
  assign sq_last = 1'b1;
  assign sq_msg = {rdma_base_params,{rdma_base_len,{rdma_base_rvaddr,rdma_base_lvaddr}}};
  assign sq_rsrvd = 14'h0;
  assign io_rdma_sq_payload_data = {sq_opcode,{sq_qpn,{sq_host,{sq_mode,{sq_last,{sq_msg,sq_rsrvd}}}}}};
  assign streamFifo_10_io_flush = (! io_ctrl_en);
  assign streamFifo_11_io_flush = (! io_ctrl_en);
  assign timeOutInc = (10'h0 < streamFifo_10_io_occupancy);
  assign io_q_sink_ready = streamFifo_10_io_push_ready;
  assign _zz_io_rdma_axis_src_valid = (8'h0 < _zz_io_rdma_sq_valid);
  assign streamFifo_10_io_pop_ready = (io_rdma_axis_src_ready && _zz_io_rdma_axis_src_valid);
  assign io_rdma_axis_src_valid = (streamFifo_10_io_pop_valid && _zz_io_rdma_axis_src_valid);
  assign io_rdma_axis_src_payload_tdata = streamFifo_10_io_pop_payload;
  assign io_rdma_sq_valid = (($signed(_zz_io_rdma_sq_valid_5) <= $signed(_zz_io_rdma_sq_valid_6)) || _zz_io_rdma_sq_valid_4);
  assign io_q_src_valid = streamFifo_11_io_pop_valid;
  assign io_q_src_payload = streamFifo_11_io_pop_payload;
  assign io_rdma_axis_sink_ready = streamFifo_11_io_push_ready;
  assign when_RdmaFlowBpss_l117 = (! io_ctrl_en);
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_rdma_sq_valid <= 8'h0;
      _zz_io_rdma_sq_valid_3 <= 9'h0;
      _zz_when_RdmaFlowBpss_l47 <= 26'h0;
    end else begin
      if((switch_Utils_l16 == {1'b1,1'b0})) begin
          _zz_io_rdma_sq_valid <= (_zz_io_rdma_sq_valid + 8'h01);
      end else if((switch_Utils_l16 == {1'b0,1'b1})) begin
          _zz_io_rdma_sq_valid <= (_zz_io_rdma_sq_valid - 8'h01);
      end
      if(when_Utils_l21) begin
        _zz_io_rdma_sq_valid <= 8'h0;
      end
      _zz_io_rdma_sq_valid_3 <= _zz_io_rdma_sq_valid_2;
      if((switch_Utils_l34 == {1'b1,1'b0})) begin
          _zz_when_RdmaFlowBpss_l47 <= (_zz_when_RdmaFlowBpss_l47 + 26'h0000001);
      end else if((switch_Utils_l34 == {1'b0,1'b1})) begin
          _zz_when_RdmaFlowBpss_l47 <= (_zz_when_RdmaFlowBpss_l47 - 26'h0000001);
      end
      if(when_Utils_l39) begin
        _zz_when_RdmaFlowBpss_l47 <= 26'h0;
      end
    end
  end

  always @(posedge clk) begin
    if(when_Utils_l63) begin
      _zz_when_Utils_l65 <= 1'b1;
    end
    if(io_rdma_sq_fire) begin
      _zz_when_Utils_l65 <= 1'b0;
    end
    if(when_RdmaFlowBpss_l44) begin
      rTimeOut <= _zz_io_rdma_sq_valid_4;
    end
  end


endmodule

module WrapNode (
  output              io_axi_0_aw_valid,
  input               io_axi_0_aw_ready,
  output     [63:0]   io_axi_0_aw_payload_addr,
  output     [5:0]    io_axi_0_aw_payload_id,
  output     [7:0]    io_axi_0_aw_payload_len,
  output     [2:0]    io_axi_0_aw_payload_size,
  output     [1:0]    io_axi_0_aw_payload_burst,
  output              io_axi_0_w_valid,
  input               io_axi_0_w_ready,
  output     [511:0]  io_axi_0_w_payload_data,
  output     [63:0]   io_axi_0_w_payload_strb,
  output              io_axi_0_w_payload_last,
  input               io_axi_0_b_valid,
  output              io_axi_0_b_ready,
  input      [5:0]    io_axi_0_b_payload_id,
  input      [1:0]    io_axi_0_b_payload_resp,
  output              io_axi_0_ar_valid,
  input               io_axi_0_ar_ready,
  output     [63:0]   io_axi_0_ar_payload_addr,
  output     [5:0]    io_axi_0_ar_payload_id,
  output     [7:0]    io_axi_0_ar_payload_len,
  output     [2:0]    io_axi_0_ar_payload_size,
  output     [1:0]    io_axi_0_ar_payload_burst,
  input               io_axi_0_r_valid,
  output              io_axi_0_r_ready,
  input      [511:0]  io_axi_0_r_payload_data,
  input      [5:0]    io_axi_0_r_payload_id,
  input      [1:0]    io_axi_0_r_payload_resp,
  input               io_axi_0_r_payload_last,
  output              io_axi_1_aw_valid,
  input               io_axi_1_aw_ready,
  output     [63:0]   io_axi_1_aw_payload_addr,
  output     [5:0]    io_axi_1_aw_payload_id,
  output     [7:0]    io_axi_1_aw_payload_len,
  output     [2:0]    io_axi_1_aw_payload_size,
  output     [1:0]    io_axi_1_aw_payload_burst,
  output              io_axi_1_w_valid,
  input               io_axi_1_w_ready,
  output     [511:0]  io_axi_1_w_payload_data,
  output     [63:0]   io_axi_1_w_payload_strb,
  output              io_axi_1_w_payload_last,
  input               io_axi_1_b_valid,
  output              io_axi_1_b_ready,
  input      [5:0]    io_axi_1_b_payload_id,
  input      [1:0]    io_axi_1_b_payload_resp,
  output              io_axi_1_ar_valid,
  input               io_axi_1_ar_ready,
  output     [63:0]   io_axi_1_ar_payload_addr,
  output     [5:0]    io_axi_1_ar_payload_id,
  output     [7:0]    io_axi_1_ar_payload_len,
  output     [2:0]    io_axi_1_ar_payload_size,
  output     [1:0]    io_axi_1_ar_payload_burst,
  input               io_axi_1_r_valid,
  output              io_axi_1_r_ready,
  input      [511:0]  io_axi_1_r_payload_data,
  input      [5:0]    io_axi_1_r_payload_id,
  input      [1:0]    io_axi_1_r_payload_resp,
  input               io_axi_1_r_payload_last,
  output              io_cmdAxi_0_aw_valid,
  input               io_cmdAxi_0_aw_ready,
  output     [63:0]   io_cmdAxi_0_aw_payload_addr,
  output     [5:0]    io_cmdAxi_0_aw_payload_id,
  output     [7:0]    io_cmdAxi_0_aw_payload_len,
  output     [2:0]    io_cmdAxi_0_aw_payload_size,
  output     [1:0]    io_cmdAxi_0_aw_payload_burst,
  output              io_cmdAxi_0_w_valid,
  input               io_cmdAxi_0_w_ready,
  output     [511:0]  io_cmdAxi_0_w_payload_data,
  output     [63:0]   io_cmdAxi_0_w_payload_strb,
  output              io_cmdAxi_0_w_payload_last,
  input               io_cmdAxi_0_b_valid,
  output              io_cmdAxi_0_b_ready,
  input      [5:0]    io_cmdAxi_0_b_payload_id,
  input      [1:0]    io_cmdAxi_0_b_payload_resp,
  output              io_cmdAxi_0_ar_valid,
  input               io_cmdAxi_0_ar_ready,
  output     [63:0]   io_cmdAxi_0_ar_payload_addr,
  output     [5:0]    io_cmdAxi_0_ar_payload_id,
  output     [7:0]    io_cmdAxi_0_ar_payload_len,
  output     [2:0]    io_cmdAxi_0_ar_payload_size,
  output     [1:0]    io_cmdAxi_0_ar_payload_burst,
  input               io_cmdAxi_0_r_valid,
  output              io_cmdAxi_0_r_ready,
  input      [511:0]  io_cmdAxi_0_r_payload_data,
  input      [5:0]    io_cmdAxi_0_r_payload_id,
  input      [1:0]    io_cmdAxi_0_r_payload_resp,
  input               io_cmdAxi_0_r_payload_last,
  input      [0:0]    io_nodeId,
  input      [31:0]   io_txnNumTotal,
  input      [31:0]   io_cmdAddrOffs_0,
  input               io_start,
  output              io_done_0,
  output     [31:0]   io_cntTxnCmt_0,
  output     [31:0]   io_cntTxnAbt_0,
  output     [31:0]   io_cntTxnLd_0,
  output     [31:0]   io_cntLockLoc_0,
  output     [31:0]   io_cntLockRmt_0,
  output     [31:0]   io_cntLockDenyLoc_0,
  output     [31:0]   io_cntLockDenyRmt_0,
  output     [31:0]   io_cntClk_0,
  output              io_sendQ_valid,
  input               io_sendQ_ready,
  output     [511:0]  io_sendQ_payload,
  output              io_respQ_valid,
  input               io_respQ_ready,
  output     [511:0]  io_respQ_payload,
  input               io_reqQ_valid,
  output              io_reqQ_ready,
  input      [511:0]  io_reqQ_payload,
  input               io_recvQ_valid,
  output              io_recvQ_ready,
  input      [511:0]  io_recvQ_payload,
  output              io_sendStatusVld,
  output              io_recvStatusVld,
  output     [3:0]    io_nReq,
  output     [3:0]    io_nWrCmtReq,
  output     [3:0]    io_nRdGetReq,
  output     [3:0]    io_nResp,
  output     [3:0]    io_nWrCmtResp,
  output     [3:0]    io_nRdGetResp,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                txnManAry_0_io_lkReqLoc_ready;
  wire                ltMCh_io_lt_0_lkResp_ready;
  wire                txnManAry_0_io_lkReqLoc_valid;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_payload_nId;
  wire       [21:0]   txnManAry_0_io_lkReqLoc_payload_tId;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_payload_tabId;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_payload_snId;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_payload_txnId;
  wire       [1:0]    txnManAry_0_io_lkReqLoc_payload_lkType;
  wire                txnManAry_0_io_lkReqLoc_payload_lkRelease;
  wire                txnManAry_0_io_lkReqLoc_payload_txnTimeOut;
  wire                txnManAry_0_io_lkReqLoc_payload_txnAbt;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_payload_lkIdx;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_payload_wLen;
  wire                txnManAry_0_io_lkReqRmt_valid;
  wire       [0:0]    txnManAry_0_io_lkReqRmt_payload_nId;
  wire       [21:0]   txnManAry_0_io_lkReqRmt_payload_tId;
  wire       [2:0]    txnManAry_0_io_lkReqRmt_payload_tabId;
  wire       [0:0]    txnManAry_0_io_lkReqRmt_payload_snId;
  wire       [5:0]    txnManAry_0_io_lkReqRmt_payload_txnId;
  wire       [1:0]    txnManAry_0_io_lkReqRmt_payload_lkType;
  wire                txnManAry_0_io_lkReqRmt_payload_lkRelease;
  wire                txnManAry_0_io_lkReqRmt_payload_txnTimeOut;
  wire                txnManAry_0_io_lkReqRmt_payload_txnAbt;
  wire       [5:0]    txnManAry_0_io_lkReqRmt_payload_lkIdx;
  wire       [2:0]    txnManAry_0_io_lkReqRmt_payload_wLen;
  wire                txnManAry_0_io_lkRespLoc_ready;
  wire                txnManAry_0_io_lkRespRmt_ready;
  wire                txnManAry_0_io_rdRmt_ready;
  wire                txnManAry_0_io_wrRmt_valid;
  wire       [511:0]  txnManAry_0_io_wrRmt_payload;
  wire                txnManAry_0_io_axi_ar_valid;
  wire       [63:0]   txnManAry_0_io_axi_ar_payload_addr;
  wire       [5:0]    txnManAry_0_io_axi_ar_payload_id;
  wire       [7:0]    txnManAry_0_io_axi_ar_payload_len;
  wire       [2:0]    txnManAry_0_io_axi_ar_payload_size;
  wire       [1:0]    txnManAry_0_io_axi_ar_payload_burst;
  wire                txnManAry_0_io_axi_aw_valid;
  wire       [63:0]   txnManAry_0_io_axi_aw_payload_addr;
  wire       [5:0]    txnManAry_0_io_axi_aw_payload_id;
  wire       [7:0]    txnManAry_0_io_axi_aw_payload_len;
  wire       [2:0]    txnManAry_0_io_axi_aw_payload_size;
  wire       [1:0]    txnManAry_0_io_axi_aw_payload_burst;
  wire                txnManAry_0_io_axi_w_valid;
  wire       [511:0]  txnManAry_0_io_axi_w_payload_data;
  wire       [63:0]   txnManAry_0_io_axi_w_payload_strb;
  wire                txnManAry_0_io_axi_w_payload_last;
  wire                txnManAry_0_io_axi_r_ready;
  wire                txnManAry_0_io_axi_b_ready;
  wire                txnManAry_0_io_cmdAxi_ar_valid;
  wire       [63:0]   txnManAry_0_io_cmdAxi_ar_payload_addr;
  wire       [5:0]    txnManAry_0_io_cmdAxi_ar_payload_id;
  wire       [7:0]    txnManAry_0_io_cmdAxi_ar_payload_len;
  wire       [2:0]    txnManAry_0_io_cmdAxi_ar_payload_size;
  wire       [1:0]    txnManAry_0_io_cmdAxi_ar_payload_burst;
  wire                txnManAry_0_io_cmdAxi_aw_valid;
  wire       [63:0]   txnManAry_0_io_cmdAxi_aw_payload_addr;
  wire       [5:0]    txnManAry_0_io_cmdAxi_aw_payload_id;
  wire       [7:0]    txnManAry_0_io_cmdAxi_aw_payload_len;
  wire       [2:0]    txnManAry_0_io_cmdAxi_aw_payload_size;
  wire       [1:0]    txnManAry_0_io_cmdAxi_aw_payload_burst;
  wire                txnManAry_0_io_cmdAxi_w_valid;
  wire       [511:0]  txnManAry_0_io_cmdAxi_w_payload_data;
  wire       [63:0]   txnManAry_0_io_cmdAxi_w_payload_strb;
  wire                txnManAry_0_io_cmdAxi_w_payload_last;
  wire                txnManAry_0_io_cmdAxi_r_ready;
  wire                txnManAry_0_io_cmdAxi_b_ready;
  wire                txnManAry_0_io_done;
  wire       [31:0]   txnManAry_0_io_cntTxnCmt;
  wire       [31:0]   txnManAry_0_io_cntTxnAbt;
  wire       [31:0]   txnManAry_0_io_cntTxnLd;
  wire       [31:0]   txnManAry_0_io_cntLockLoc;
  wire       [31:0]   txnManAry_0_io_cntLockRmt;
  wire       [31:0]   txnManAry_0_io_cntLockDenyLoc;
  wire       [31:0]   txnManAry_0_io_cntLockDenyRmt;
  wire       [31:0]   txnManAry_0_io_cntClk;
  wire                ltMCh_io_lt_0_lkReq_ready;
  wire                ltMCh_io_lt_0_lkResp_valid;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_payload_nId;
  wire       [21:0]   ltMCh_io_lt_0_lkResp_payload_tId;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_payload_tabId;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_payload_snId;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_payload_txnId;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_payload_lkType;
  wire                ltMCh_io_lt_0_lkResp_payload_lkRelease;
  wire                ltMCh_io_lt_0_lkResp_payload_txnAbt;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_payload_lkIdx;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_payload_wLen;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_payload_respType;
  wire                ltMCh_io_lt_0_lkResp_payload_lkWaited;
  wire                ltMCh_io_lt_1_lkReq_ready;
  wire                ltMCh_io_lt_1_lkResp_valid;
  wire       [0:0]    ltMCh_io_lt_1_lkResp_payload_nId;
  wire       [21:0]   ltMCh_io_lt_1_lkResp_payload_tId;
  wire       [2:0]    ltMCh_io_lt_1_lkResp_payload_tabId;
  wire       [0:0]    ltMCh_io_lt_1_lkResp_payload_snId;
  wire       [5:0]    ltMCh_io_lt_1_lkResp_payload_txnId;
  wire       [1:0]    ltMCh_io_lt_1_lkResp_payload_lkType;
  wire                ltMCh_io_lt_1_lkResp_payload_lkRelease;
  wire                ltMCh_io_lt_1_lkResp_payload_txnAbt;
  wire       [5:0]    ltMCh_io_lt_1_lkResp_payload_lkIdx;
  wire       [2:0]    ltMCh_io_lt_1_lkResp_payload_wLen;
  wire       [1:0]    ltMCh_io_lt_1_lkResp_payload_respType;
  wire                ltMCh_io_lt_1_lkResp_payload_lkWaited;
  wire                txnAgent_1_io_lkReq_ready;
  wire                txnAgent_1_io_wrData_ready;
  wire                txnAgent_1_io_lkResp_valid;
  wire       [0:0]    txnAgent_1_io_lkResp_payload_nId;
  wire       [21:0]   txnAgent_1_io_lkResp_payload_tId;
  wire       [2:0]    txnAgent_1_io_lkResp_payload_tabId;
  wire       [0:0]    txnAgent_1_io_lkResp_payload_snId;
  wire       [5:0]    txnAgent_1_io_lkResp_payload_txnId;
  wire       [1:0]    txnAgent_1_io_lkResp_payload_lkType;
  wire                txnAgent_1_io_lkResp_payload_lkRelease;
  wire                txnAgent_1_io_lkResp_payload_txnAbt;
  wire       [5:0]    txnAgent_1_io_lkResp_payload_lkIdx;
  wire       [2:0]    txnAgent_1_io_lkResp_payload_wLen;
  wire       [1:0]    txnAgent_1_io_lkResp_payload_respType;
  wire                txnAgent_1_io_lkResp_payload_lkWaited;
  wire                txnAgent_1_io_rdData_valid;
  wire       [511:0]  txnAgent_1_io_rdData_payload;
  wire                txnAgent_1_io_axi_ar_valid;
  wire       [63:0]   txnAgent_1_io_axi_ar_payload_addr;
  wire       [5:0]    txnAgent_1_io_axi_ar_payload_id;
  wire       [7:0]    txnAgent_1_io_axi_ar_payload_len;
  wire       [2:0]    txnAgent_1_io_axi_ar_payload_size;
  wire       [1:0]    txnAgent_1_io_axi_ar_payload_burst;
  wire                txnAgent_1_io_axi_aw_valid;
  wire       [63:0]   txnAgent_1_io_axi_aw_payload_addr;
  wire       [5:0]    txnAgent_1_io_axi_aw_payload_id;
  wire       [7:0]    txnAgent_1_io_axi_aw_payload_len;
  wire       [2:0]    txnAgent_1_io_axi_aw_payload_size;
  wire       [1:0]    txnAgent_1_io_axi_aw_payload_burst;
  wire                txnAgent_1_io_axi_w_valid;
  wire       [511:0]  txnAgent_1_io_axi_w_payload_data;
  wire       [63:0]   txnAgent_1_io_axi_w_payload_strb;
  wire                txnAgent_1_io_axi_w_payload_last;
  wire                txnAgent_1_io_axi_r_ready;
  wire                txnAgent_1_io_axi_b_ready;
  wire                txnAgent_1_io_ltReq_valid;
  wire       [0:0]    txnAgent_1_io_ltReq_payload_nId;
  wire       [21:0]   txnAgent_1_io_ltReq_payload_tId;
  wire       [2:0]    txnAgent_1_io_ltReq_payload_tabId;
  wire       [0:0]    txnAgent_1_io_ltReq_payload_snId;
  wire       [5:0]    txnAgent_1_io_ltReq_payload_txnId;
  wire       [1:0]    txnAgent_1_io_ltReq_payload_lkType;
  wire                txnAgent_1_io_ltReq_payload_lkRelease;
  wire                txnAgent_1_io_ltReq_payload_txnTimeOut;
  wire                txnAgent_1_io_ltReq_payload_txnAbt;
  wire       [5:0]    txnAgent_1_io_ltReq_payload_lkIdx;
  wire       [2:0]    txnAgent_1_io_ltReq_payload_wLen;
  wire                txnAgent_1_io_ltResp_ready;
  wire                sendArb_io_lkReqV_0_ready;
  wire                sendArb_io_wrDataV_0_ready;
  wire                sendArb_io_sendQ_valid;
  wire       [511:0]  sendArb_io_sendQ_payload;
  wire                sendArb_io_statusVld;
  wire       [3:0]    sendArb_io_nReq;
  wire       [3:0]    sendArb_io_nWrCmtReq;
  wire       [3:0]    sendArb_io_nRdGetReq;
  wire                recvDisp_io_recvQ_ready;
  wire                recvDisp_io_lkRespV_0_valid;
  wire       [0:0]    recvDisp_io_lkRespV_0_payload_nId;
  wire       [21:0]   recvDisp_io_lkRespV_0_payload_tId;
  wire       [2:0]    recvDisp_io_lkRespV_0_payload_tabId;
  wire       [0:0]    recvDisp_io_lkRespV_0_payload_snId;
  wire       [5:0]    recvDisp_io_lkRespV_0_payload_txnId;
  wire       [1:0]    recvDisp_io_lkRespV_0_payload_lkType;
  wire                recvDisp_io_lkRespV_0_payload_lkRelease;
  wire                recvDisp_io_lkRespV_0_payload_txnAbt;
  wire       [5:0]    recvDisp_io_lkRespV_0_payload_lkIdx;
  wire       [2:0]    recvDisp_io_lkRespV_0_payload_wLen;
  wire       [1:0]    recvDisp_io_lkRespV_0_payload_respType;
  wire                recvDisp_io_lkRespV_0_payload_lkWaited;
  wire                recvDisp_io_rdDataV_0_valid;
  wire       [511:0]  recvDisp_io_rdDataV_0_payload;
  wire                recvDisp_io_statusVld;
  wire       [3:0]    recvDisp_io_nResp;
  wire       [3:0]    recvDisp_io_nWrCmtResp;
  wire       [3:0]    recvDisp_io_nRdGetResp;
  wire                reqDisp_io_reqQ_ready;
  wire                reqDisp_io_lkReq_valid;
  wire       [0:0]    reqDisp_io_lkReq_payload_nId;
  wire       [21:0]   reqDisp_io_lkReq_payload_tId;
  wire       [2:0]    reqDisp_io_lkReq_payload_tabId;
  wire       [0:0]    reqDisp_io_lkReq_payload_snId;
  wire       [5:0]    reqDisp_io_lkReq_payload_txnId;
  wire       [1:0]    reqDisp_io_lkReq_payload_lkType;
  wire                reqDisp_io_lkReq_payload_lkRelease;
  wire                reqDisp_io_lkReq_payload_txnTimeOut;
  wire                reqDisp_io_lkReq_payload_txnAbt;
  wire       [5:0]    reqDisp_io_lkReq_payload_lkIdx;
  wire       [2:0]    reqDisp_io_lkReq_payload_wLen;
  wire                reqDisp_io_wrData_valid;
  wire       [511:0]  reqDisp_io_wrData_payload;
  wire                respArb_io_lkResp_ready;
  wire                respArb_io_rdData_ready;
  wire                respArb_io_respQ_valid;
  wire       [511:0]  respArb_io_respQ_payload;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_valid;
  reg                 txnManAry_0_io_lkReqLoc_s2mPipe_ready;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_nId;
  wire       [21:0]   txnManAry_0_io_lkReqLoc_s2mPipe_payload_tId;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_tabId;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_snId;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnId;
  wire       [1:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkRelease;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnTimeOut;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnAbt;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkIdx;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_payload_wLen;
  reg                 txnManAry_0_io_lkReqLoc_rValid;
  reg        [0:0]    txnManAry_0_io_lkReqLoc_rData_nId;
  reg        [21:0]   txnManAry_0_io_lkReqLoc_rData_tId;
  reg        [2:0]    txnManAry_0_io_lkReqLoc_rData_tabId;
  reg        [0:0]    txnManAry_0_io_lkReqLoc_rData_snId;
  reg        [5:0]    txnManAry_0_io_lkReqLoc_rData_txnId;
  reg        [1:0]    txnManAry_0_io_lkReqLoc_rData_lkType;
  reg                 txnManAry_0_io_lkReqLoc_rData_lkRelease;
  reg                 txnManAry_0_io_lkReqLoc_rData_txnTimeOut;
  reg                 txnManAry_0_io_lkReqLoc_rData_txnAbt;
  reg        [5:0]    txnManAry_0_io_lkReqLoc_rData_lkIdx;
  reg        [2:0]    txnManAry_0_io_lkReqLoc_rData_wLen;
  wire       [1:0]    _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_valid;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_ready;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkRelease;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_wLen;
  reg                 txnManAry_0_io_lkReqLoc_s2mPipe_rValid;
  reg        [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_nId;
  reg        [21:0]   txnManAry_0_io_lkReqLoc_s2mPipe_rData_tId;
  reg        [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_tabId;
  reg        [0:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_snId;
  reg        [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnId;
  reg        [1:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType;
  reg                 txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkRelease;
  reg                 txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnTimeOut;
  reg                 txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnAbt;
  reg        [5:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkIdx;
  reg        [2:0]    txnManAry_0_io_lkReqLoc_s2mPipe_rData_wLen;
  wire                when_Stream_l368;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_valid;
  reg                 ltMCh_io_lt_0_lkResp_s2mPipe_ready;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_nId;
  wire       [21:0]   ltMCh_io_lt_0_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkRelease;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltMCh_io_lt_0_lkResp_rValid;
  reg        [0:0]    ltMCh_io_lt_0_lkResp_rData_nId;
  reg        [21:0]   ltMCh_io_lt_0_lkResp_rData_tId;
  reg        [2:0]    ltMCh_io_lt_0_lkResp_rData_tabId;
  reg        [0:0]    ltMCh_io_lt_0_lkResp_rData_snId;
  reg        [5:0]    ltMCh_io_lt_0_lkResp_rData_txnId;
  reg        [1:0]    ltMCh_io_lt_0_lkResp_rData_lkType;
  reg                 ltMCh_io_lt_0_lkResp_rData_lkRelease;
  reg                 ltMCh_io_lt_0_lkResp_rData_txnAbt;
  reg        [5:0]    ltMCh_io_lt_0_lkResp_rData_lkIdx;
  reg        [2:0]    ltMCh_io_lt_0_lkResp_rData_wLen;
  reg        [1:0]    ltMCh_io_lt_0_lkResp_rData_respType;
  reg                 ltMCh_io_lt_0_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltMCh_io_lt_0_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_nId;
  reg        [21:0]   ltMCh_io_lt_0_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType;
  reg                 ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType;
  reg                 ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_1;
  `ifndef SYNTHESIS
  reg [47:0] txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string;
  reg [47:0] txnManAry_0_io_lkReqLoc_rData_lkType_string;
  reg [47:0] _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string;
  reg [47:0] txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string;
  reg [47:0] ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltMCh_io_lt_0_lkResp_rData_lkType_string;
  reg [71:0] ltMCh_io_lt_0_lkResp_rData_respType_string;
  reg [47:0] _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string;
  `endif


  TxnManCS txnManAry_0 (
    .io_lkReqLoc_valid              (txnManAry_0_io_lkReqLoc_valid                             ), //o
    .io_lkReqLoc_ready              (txnManAry_0_io_lkReqLoc_ready                             ), //i
    .io_lkReqLoc_payload_nId        (txnManAry_0_io_lkReqLoc_payload_nId                       ), //o
    .io_lkReqLoc_payload_tId        (txnManAry_0_io_lkReqLoc_payload_tId[21:0]                 ), //o
    .io_lkReqLoc_payload_tabId      (txnManAry_0_io_lkReqLoc_payload_tabId[2:0]                ), //o
    .io_lkReqLoc_payload_snId       (txnManAry_0_io_lkReqLoc_payload_snId                      ), //o
    .io_lkReqLoc_payload_txnId      (txnManAry_0_io_lkReqLoc_payload_txnId[5:0]                ), //o
    .io_lkReqLoc_payload_lkType     (txnManAry_0_io_lkReqLoc_payload_lkType[1:0]               ), //o
    .io_lkReqLoc_payload_lkRelease  (txnManAry_0_io_lkReqLoc_payload_lkRelease                 ), //o
    .io_lkReqLoc_payload_txnTimeOut (txnManAry_0_io_lkReqLoc_payload_txnTimeOut                ), //o
    .io_lkReqLoc_payload_txnAbt     (txnManAry_0_io_lkReqLoc_payload_txnAbt                    ), //o
    .io_lkReqLoc_payload_lkIdx      (txnManAry_0_io_lkReqLoc_payload_lkIdx[5:0]                ), //o
    .io_lkReqLoc_payload_wLen       (txnManAry_0_io_lkReqLoc_payload_wLen[2:0]                 ), //o
    .io_lkReqRmt_valid              (txnManAry_0_io_lkReqRmt_valid                             ), //o
    .io_lkReqRmt_ready              (sendArb_io_lkReqV_0_ready                                 ), //i
    .io_lkReqRmt_payload_nId        (txnManAry_0_io_lkReqRmt_payload_nId                       ), //o
    .io_lkReqRmt_payload_tId        (txnManAry_0_io_lkReqRmt_payload_tId[21:0]                 ), //o
    .io_lkReqRmt_payload_tabId      (txnManAry_0_io_lkReqRmt_payload_tabId[2:0]                ), //o
    .io_lkReqRmt_payload_snId       (txnManAry_0_io_lkReqRmt_payload_snId                      ), //o
    .io_lkReqRmt_payload_txnId      (txnManAry_0_io_lkReqRmt_payload_txnId[5:0]                ), //o
    .io_lkReqRmt_payload_lkType     (txnManAry_0_io_lkReqRmt_payload_lkType[1:0]               ), //o
    .io_lkReqRmt_payload_lkRelease  (txnManAry_0_io_lkReqRmt_payload_lkRelease                 ), //o
    .io_lkReqRmt_payload_txnTimeOut (txnManAry_0_io_lkReqRmt_payload_txnTimeOut                ), //o
    .io_lkReqRmt_payload_txnAbt     (txnManAry_0_io_lkReqRmt_payload_txnAbt                    ), //o
    .io_lkReqRmt_payload_lkIdx      (txnManAry_0_io_lkReqRmt_payload_lkIdx[5:0]                ), //o
    .io_lkReqRmt_payload_wLen       (txnManAry_0_io_lkReqRmt_payload_wLen[2:0]                 ), //o
    .io_lkRespLoc_valid             (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_lkRespLoc_ready             (txnManAry_0_io_lkRespLoc_ready                            ), //o
    .io_lkRespLoc_payload_nId       (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_lkRespLoc_payload_tId       (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tId[21:0]    ), //i
    .io_lkRespLoc_payload_tabId     (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_lkRespLoc_payload_snId      (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_lkRespLoc_payload_txnId     (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_lkRespLoc_payload_lkType    (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_lkRespLoc_payload_lkRelease (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_lkRespLoc_payload_txnAbt    (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_lkRespLoc_payload_lkIdx     (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_lkRespLoc_payload_wLen      (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_lkRespLoc_payload_respType  (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_lkRespLoc_payload_lkWaited  (ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_lkRespRmt_valid             (recvDisp_io_lkRespV_0_valid                               ), //i
    .io_lkRespRmt_ready             (txnManAry_0_io_lkRespRmt_ready                            ), //o
    .io_lkRespRmt_payload_nId       (recvDisp_io_lkRespV_0_payload_nId                         ), //i
    .io_lkRespRmt_payload_tId       (recvDisp_io_lkRespV_0_payload_tId[21:0]                   ), //i
    .io_lkRespRmt_payload_tabId     (recvDisp_io_lkRespV_0_payload_tabId[2:0]                  ), //i
    .io_lkRespRmt_payload_snId      (recvDisp_io_lkRespV_0_payload_snId                        ), //i
    .io_lkRespRmt_payload_txnId     (recvDisp_io_lkRespV_0_payload_txnId[5:0]                  ), //i
    .io_lkRespRmt_payload_lkType    (recvDisp_io_lkRespV_0_payload_lkType[1:0]                 ), //i
    .io_lkRespRmt_payload_lkRelease (recvDisp_io_lkRespV_0_payload_lkRelease                   ), //i
    .io_lkRespRmt_payload_txnAbt    (recvDisp_io_lkRespV_0_payload_txnAbt                      ), //i
    .io_lkRespRmt_payload_lkIdx     (recvDisp_io_lkRespV_0_payload_lkIdx[5:0]                  ), //i
    .io_lkRespRmt_payload_wLen      (recvDisp_io_lkRespV_0_payload_wLen[2:0]                   ), //i
    .io_lkRespRmt_payload_respType  (recvDisp_io_lkRespV_0_payload_respType[1:0]               ), //i
    .io_lkRespRmt_payload_lkWaited  (recvDisp_io_lkRespV_0_payload_lkWaited                    ), //i
    .io_rdRmt_valid                 (recvDisp_io_rdDataV_0_valid                               ), //i
    .io_rdRmt_ready                 (txnManAry_0_io_rdRmt_ready                                ), //o
    .io_rdRmt_payload               (recvDisp_io_rdDataV_0_payload[511:0]                      ), //i
    .io_wrRmt_valid                 (txnManAry_0_io_wrRmt_valid                                ), //o
    .io_wrRmt_ready                 (sendArb_io_wrDataV_0_ready                                ), //i
    .io_wrRmt_payload               (txnManAry_0_io_wrRmt_payload[511:0]                       ), //o
    .io_axi_aw_valid                (txnManAry_0_io_axi_aw_valid                               ), //o
    .io_axi_aw_ready                (io_axi_0_aw_ready                                         ), //i
    .io_axi_aw_payload_addr         (txnManAry_0_io_axi_aw_payload_addr[63:0]                  ), //o
    .io_axi_aw_payload_id           (txnManAry_0_io_axi_aw_payload_id[5:0]                     ), //o
    .io_axi_aw_payload_len          (txnManAry_0_io_axi_aw_payload_len[7:0]                    ), //o
    .io_axi_aw_payload_size         (txnManAry_0_io_axi_aw_payload_size[2:0]                   ), //o
    .io_axi_aw_payload_burst        (txnManAry_0_io_axi_aw_payload_burst[1:0]                  ), //o
    .io_axi_w_valid                 (txnManAry_0_io_axi_w_valid                                ), //o
    .io_axi_w_ready                 (io_axi_0_w_ready                                          ), //i
    .io_axi_w_payload_data          (txnManAry_0_io_axi_w_payload_data[511:0]                  ), //o
    .io_axi_w_payload_strb          (txnManAry_0_io_axi_w_payload_strb[63:0]                   ), //o
    .io_axi_w_payload_last          (txnManAry_0_io_axi_w_payload_last                         ), //o
    .io_axi_b_valid                 (io_axi_0_b_valid                                          ), //i
    .io_axi_b_ready                 (txnManAry_0_io_axi_b_ready                                ), //o
    .io_axi_b_payload_id            (io_axi_0_b_payload_id[5:0]                                ), //i
    .io_axi_b_payload_resp          (io_axi_0_b_payload_resp[1:0]                              ), //i
    .io_axi_ar_valid                (txnManAry_0_io_axi_ar_valid                               ), //o
    .io_axi_ar_ready                (io_axi_0_ar_ready                                         ), //i
    .io_axi_ar_payload_addr         (txnManAry_0_io_axi_ar_payload_addr[63:0]                  ), //o
    .io_axi_ar_payload_id           (txnManAry_0_io_axi_ar_payload_id[5:0]                     ), //o
    .io_axi_ar_payload_len          (txnManAry_0_io_axi_ar_payload_len[7:0]                    ), //o
    .io_axi_ar_payload_size         (txnManAry_0_io_axi_ar_payload_size[2:0]                   ), //o
    .io_axi_ar_payload_burst        (txnManAry_0_io_axi_ar_payload_burst[1:0]                  ), //o
    .io_axi_r_valid                 (io_axi_0_r_valid                                          ), //i
    .io_axi_r_ready                 (txnManAry_0_io_axi_r_ready                                ), //o
    .io_axi_r_payload_data          (io_axi_0_r_payload_data[511:0]                            ), //i
    .io_axi_r_payload_id            (io_axi_0_r_payload_id[5:0]                                ), //i
    .io_axi_r_payload_resp          (io_axi_0_r_payload_resp[1:0]                              ), //i
    .io_axi_r_payload_last          (io_axi_0_r_payload_last                                   ), //i
    .io_cmdAxi_aw_valid             (txnManAry_0_io_cmdAxi_aw_valid                            ), //o
    .io_cmdAxi_aw_ready             (io_cmdAxi_0_aw_ready                                      ), //i
    .io_cmdAxi_aw_payload_addr      (txnManAry_0_io_cmdAxi_aw_payload_addr[63:0]               ), //o
    .io_cmdAxi_aw_payload_id        (txnManAry_0_io_cmdAxi_aw_payload_id[5:0]                  ), //o
    .io_cmdAxi_aw_payload_len       (txnManAry_0_io_cmdAxi_aw_payload_len[7:0]                 ), //o
    .io_cmdAxi_aw_payload_size      (txnManAry_0_io_cmdAxi_aw_payload_size[2:0]                ), //o
    .io_cmdAxi_aw_payload_burst     (txnManAry_0_io_cmdAxi_aw_payload_burst[1:0]               ), //o
    .io_cmdAxi_w_valid              (txnManAry_0_io_cmdAxi_w_valid                             ), //o
    .io_cmdAxi_w_ready              (io_cmdAxi_0_w_ready                                       ), //i
    .io_cmdAxi_w_payload_data       (txnManAry_0_io_cmdAxi_w_payload_data[511:0]               ), //o
    .io_cmdAxi_w_payload_strb       (txnManAry_0_io_cmdAxi_w_payload_strb[63:0]                ), //o
    .io_cmdAxi_w_payload_last       (txnManAry_0_io_cmdAxi_w_payload_last                      ), //o
    .io_cmdAxi_b_valid              (io_cmdAxi_0_b_valid                                       ), //i
    .io_cmdAxi_b_ready              (txnManAry_0_io_cmdAxi_b_ready                             ), //o
    .io_cmdAxi_b_payload_id         (io_cmdAxi_0_b_payload_id[5:0]                             ), //i
    .io_cmdAxi_b_payload_resp       (io_cmdAxi_0_b_payload_resp[1:0]                           ), //i
    .io_cmdAxi_ar_valid             (txnManAry_0_io_cmdAxi_ar_valid                            ), //o
    .io_cmdAxi_ar_ready             (io_cmdAxi_0_ar_ready                                      ), //i
    .io_cmdAxi_ar_payload_addr      (txnManAry_0_io_cmdAxi_ar_payload_addr[63:0]               ), //o
    .io_cmdAxi_ar_payload_id        (txnManAry_0_io_cmdAxi_ar_payload_id[5:0]                  ), //o
    .io_cmdAxi_ar_payload_len       (txnManAry_0_io_cmdAxi_ar_payload_len[7:0]                 ), //o
    .io_cmdAxi_ar_payload_size      (txnManAry_0_io_cmdAxi_ar_payload_size[2:0]                ), //o
    .io_cmdAxi_ar_payload_burst     (txnManAry_0_io_cmdAxi_ar_payload_burst[1:0]               ), //o
    .io_cmdAxi_r_valid              (io_cmdAxi_0_r_valid                                       ), //i
    .io_cmdAxi_r_ready              (txnManAry_0_io_cmdAxi_r_ready                             ), //o
    .io_cmdAxi_r_payload_data       (io_cmdAxi_0_r_payload_data[511:0]                         ), //i
    .io_cmdAxi_r_payload_id         (io_cmdAxi_0_r_payload_id[5:0]                             ), //i
    .io_cmdAxi_r_payload_resp       (io_cmdAxi_0_r_payload_resp[1:0]                           ), //i
    .io_cmdAxi_r_payload_last       (io_cmdAxi_0_r_payload_last                                ), //i
    .io_start                       (io_start                                                  ), //i
    .io_nodeId                      (io_nodeId                                                 ), //i
    .io_txnNumTotal                 (io_txnNumTotal[31:0]                                      ), //i
    .io_cmdAddrOffs                 (io_cmdAddrOffs_0[31:0]                                    ), //i
    .io_done                        (txnManAry_0_io_done                                       ), //o
    .io_cntTxnCmt                   (txnManAry_0_io_cntTxnCmt[31:0]                            ), //o
    .io_cntTxnAbt                   (txnManAry_0_io_cntTxnAbt[31:0]                            ), //o
    .io_cntTxnLd                    (txnManAry_0_io_cntTxnLd[31:0]                             ), //o
    .io_cntLockLoc                  (txnManAry_0_io_cntLockLoc[31:0]                           ), //o
    .io_cntLockRmt                  (txnManAry_0_io_cntLockRmt[31:0]                           ), //o
    .io_cntLockDenyLoc              (txnManAry_0_io_cntLockDenyLoc[31:0]                       ), //o
    .io_cntLockDenyRmt              (txnManAry_0_io_cntLockDenyRmt[31:0]                       ), //o
    .io_cntClk                      (txnManAry_0_io_cntClk[31:0]                               ), //o
    .clk                            (clk                                                       ), //i
    .resetn                         (resetn                                                    )  //i
  );
  LtTop ltMCh (
    .io_nodeId                        (io_nodeId                                                  ), //i
    .io_lt_0_lkReq_valid              (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_valid              ), //i
    .io_lt_0_lkReq_ready              (ltMCh_io_lt_0_lkReq_ready                                  ), //o
    .io_lt_0_lkReq_payload_nId        (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lt_0_lkReq_payload_tId        (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tId[21:0]  ), //i
    .io_lt_0_lkReq_payload_tabId      (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lt_0_lkReq_payload_snId       (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lt_0_lkReq_payload_txnId      (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lt_0_lkReq_payload_lkType     (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lt_0_lkReq_payload_lkRelease  (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lt_0_lkReq_payload_txnTimeOut (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lt_0_lkReq_payload_txnAbt     (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lt_0_lkReq_payload_lkIdx      (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lt_0_lkReq_payload_wLen       (txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lt_0_lkResp_valid             (ltMCh_io_lt_0_lkResp_valid                                 ), //o
    .io_lt_0_lkResp_ready             (ltMCh_io_lt_0_lkResp_ready                                 ), //i
    .io_lt_0_lkResp_payload_nId       (ltMCh_io_lt_0_lkResp_payload_nId                           ), //o
    .io_lt_0_lkResp_payload_tId       (ltMCh_io_lt_0_lkResp_payload_tId[21:0]                     ), //o
    .io_lt_0_lkResp_payload_tabId     (ltMCh_io_lt_0_lkResp_payload_tabId[2:0]                    ), //o
    .io_lt_0_lkResp_payload_snId      (ltMCh_io_lt_0_lkResp_payload_snId                          ), //o
    .io_lt_0_lkResp_payload_txnId     (ltMCh_io_lt_0_lkResp_payload_txnId[5:0]                    ), //o
    .io_lt_0_lkResp_payload_lkType    (ltMCh_io_lt_0_lkResp_payload_lkType[1:0]                   ), //o
    .io_lt_0_lkResp_payload_lkRelease (ltMCh_io_lt_0_lkResp_payload_lkRelease                     ), //o
    .io_lt_0_lkResp_payload_txnAbt    (ltMCh_io_lt_0_lkResp_payload_txnAbt                        ), //o
    .io_lt_0_lkResp_payload_lkIdx     (ltMCh_io_lt_0_lkResp_payload_lkIdx[5:0]                    ), //o
    .io_lt_0_lkResp_payload_wLen      (ltMCh_io_lt_0_lkResp_payload_wLen[2:0]                     ), //o
    .io_lt_0_lkResp_payload_respType  (ltMCh_io_lt_0_lkResp_payload_respType[1:0]                 ), //o
    .io_lt_0_lkResp_payload_lkWaited  (ltMCh_io_lt_0_lkResp_payload_lkWaited                      ), //o
    .io_lt_1_lkReq_valid              (txnAgent_1_io_ltReq_valid                                  ), //i
    .io_lt_1_lkReq_ready              (ltMCh_io_lt_1_lkReq_ready                                  ), //o
    .io_lt_1_lkReq_payload_nId        (txnAgent_1_io_ltReq_payload_nId                            ), //i
    .io_lt_1_lkReq_payload_tId        (txnAgent_1_io_ltReq_payload_tId[21:0]                      ), //i
    .io_lt_1_lkReq_payload_tabId      (txnAgent_1_io_ltReq_payload_tabId[2:0]                     ), //i
    .io_lt_1_lkReq_payload_snId       (txnAgent_1_io_ltReq_payload_snId                           ), //i
    .io_lt_1_lkReq_payload_txnId      (txnAgent_1_io_ltReq_payload_txnId[5:0]                     ), //i
    .io_lt_1_lkReq_payload_lkType     (txnAgent_1_io_ltReq_payload_lkType[1:0]                    ), //i
    .io_lt_1_lkReq_payload_lkRelease  (txnAgent_1_io_ltReq_payload_lkRelease                      ), //i
    .io_lt_1_lkReq_payload_txnTimeOut (txnAgent_1_io_ltReq_payload_txnTimeOut                     ), //i
    .io_lt_1_lkReq_payload_txnAbt     (txnAgent_1_io_ltReq_payload_txnAbt                         ), //i
    .io_lt_1_lkReq_payload_lkIdx      (txnAgent_1_io_ltReq_payload_lkIdx[5:0]                     ), //i
    .io_lt_1_lkReq_payload_wLen       (txnAgent_1_io_ltReq_payload_wLen[2:0]                      ), //i
    .io_lt_1_lkResp_valid             (ltMCh_io_lt_1_lkResp_valid                                 ), //o
    .io_lt_1_lkResp_ready             (txnAgent_1_io_ltResp_ready                                 ), //i
    .io_lt_1_lkResp_payload_nId       (ltMCh_io_lt_1_lkResp_payload_nId                           ), //o
    .io_lt_1_lkResp_payload_tId       (ltMCh_io_lt_1_lkResp_payload_tId[21:0]                     ), //o
    .io_lt_1_lkResp_payload_tabId     (ltMCh_io_lt_1_lkResp_payload_tabId[2:0]                    ), //o
    .io_lt_1_lkResp_payload_snId      (ltMCh_io_lt_1_lkResp_payload_snId                          ), //o
    .io_lt_1_lkResp_payload_txnId     (ltMCh_io_lt_1_lkResp_payload_txnId[5:0]                    ), //o
    .io_lt_1_lkResp_payload_lkType    (ltMCh_io_lt_1_lkResp_payload_lkType[1:0]                   ), //o
    .io_lt_1_lkResp_payload_lkRelease (ltMCh_io_lt_1_lkResp_payload_lkRelease                     ), //o
    .io_lt_1_lkResp_payload_txnAbt    (ltMCh_io_lt_1_lkResp_payload_txnAbt                        ), //o
    .io_lt_1_lkResp_payload_lkIdx     (ltMCh_io_lt_1_lkResp_payload_lkIdx[5:0]                    ), //o
    .io_lt_1_lkResp_payload_wLen      (ltMCh_io_lt_1_lkResp_payload_wLen[2:0]                     ), //o
    .io_lt_1_lkResp_payload_respType  (ltMCh_io_lt_1_lkResp_payload_respType[1:0]                 ), //o
    .io_lt_1_lkResp_payload_lkWaited  (ltMCh_io_lt_1_lkResp_payload_lkWaited                      ), //o
    .resetn                           (resetn                                                     ), //i
    .clk                              (clk                                                        )  //i
  );
  TxnAgent txnAgent_1 (
    .io_lkReq_valid              (reqDisp_io_lkReq_valid                    ), //i
    .io_lkReq_ready              (txnAgent_1_io_lkReq_ready                 ), //o
    .io_lkReq_payload_nId        (reqDisp_io_lkReq_payload_nId              ), //i
    .io_lkReq_payload_tId        (reqDisp_io_lkReq_payload_tId[21:0]        ), //i
    .io_lkReq_payload_tabId      (reqDisp_io_lkReq_payload_tabId[2:0]       ), //i
    .io_lkReq_payload_snId       (reqDisp_io_lkReq_payload_snId             ), //i
    .io_lkReq_payload_txnId      (reqDisp_io_lkReq_payload_txnId[5:0]       ), //i
    .io_lkReq_payload_lkType     (reqDisp_io_lkReq_payload_lkType[1:0]      ), //i
    .io_lkReq_payload_lkRelease  (reqDisp_io_lkReq_payload_lkRelease        ), //i
    .io_lkReq_payload_txnTimeOut (reqDisp_io_lkReq_payload_txnTimeOut       ), //i
    .io_lkReq_payload_txnAbt     (reqDisp_io_lkReq_payload_txnAbt           ), //i
    .io_lkReq_payload_lkIdx      (reqDisp_io_lkReq_payload_lkIdx[5:0]       ), //i
    .io_lkReq_payload_wLen       (reqDisp_io_lkReq_payload_wLen[2:0]        ), //i
    .io_wrData_valid             (reqDisp_io_wrData_valid                   ), //i
    .io_wrData_ready             (txnAgent_1_io_wrData_ready                ), //o
    .io_wrData_payload           (reqDisp_io_wrData_payload[511:0]          ), //i
    .io_lkResp_valid             (txnAgent_1_io_lkResp_valid                ), //o
    .io_lkResp_ready             (respArb_io_lkResp_ready                   ), //i
    .io_lkResp_payload_nId       (txnAgent_1_io_lkResp_payload_nId          ), //o
    .io_lkResp_payload_tId       (txnAgent_1_io_lkResp_payload_tId[21:0]    ), //o
    .io_lkResp_payload_tabId     (txnAgent_1_io_lkResp_payload_tabId[2:0]   ), //o
    .io_lkResp_payload_snId      (txnAgent_1_io_lkResp_payload_snId         ), //o
    .io_lkResp_payload_txnId     (txnAgent_1_io_lkResp_payload_txnId[5:0]   ), //o
    .io_lkResp_payload_lkType    (txnAgent_1_io_lkResp_payload_lkType[1:0]  ), //o
    .io_lkResp_payload_lkRelease (txnAgent_1_io_lkResp_payload_lkRelease    ), //o
    .io_lkResp_payload_txnAbt    (txnAgent_1_io_lkResp_payload_txnAbt       ), //o
    .io_lkResp_payload_lkIdx     (txnAgent_1_io_lkResp_payload_lkIdx[5:0]   ), //o
    .io_lkResp_payload_wLen      (txnAgent_1_io_lkResp_payload_wLen[2:0]    ), //o
    .io_lkResp_payload_respType  (txnAgent_1_io_lkResp_payload_respType[1:0]), //o
    .io_lkResp_payload_lkWaited  (txnAgent_1_io_lkResp_payload_lkWaited     ), //o
    .io_rdData_valid             (txnAgent_1_io_rdData_valid                ), //o
    .io_rdData_ready             (respArb_io_rdData_ready                   ), //i
    .io_rdData_payload           (txnAgent_1_io_rdData_payload[511:0]       ), //o
    .io_axi_aw_valid             (txnAgent_1_io_axi_aw_valid                ), //o
    .io_axi_aw_ready             (io_axi_1_aw_ready                         ), //i
    .io_axi_aw_payload_addr      (txnAgent_1_io_axi_aw_payload_addr[63:0]   ), //o
    .io_axi_aw_payload_id        (txnAgent_1_io_axi_aw_payload_id[5:0]      ), //o
    .io_axi_aw_payload_len       (txnAgent_1_io_axi_aw_payload_len[7:0]     ), //o
    .io_axi_aw_payload_size      (txnAgent_1_io_axi_aw_payload_size[2:0]    ), //o
    .io_axi_aw_payload_burst     (txnAgent_1_io_axi_aw_payload_burst[1:0]   ), //o
    .io_axi_w_valid              (txnAgent_1_io_axi_w_valid                 ), //o
    .io_axi_w_ready              (io_axi_1_w_ready                          ), //i
    .io_axi_w_payload_data       (txnAgent_1_io_axi_w_payload_data[511:0]   ), //o
    .io_axi_w_payload_strb       (txnAgent_1_io_axi_w_payload_strb[63:0]    ), //o
    .io_axi_w_payload_last       (txnAgent_1_io_axi_w_payload_last          ), //o
    .io_axi_b_valid              (io_axi_1_b_valid                          ), //i
    .io_axi_b_ready              (txnAgent_1_io_axi_b_ready                 ), //o
    .io_axi_b_payload_id         (io_axi_1_b_payload_id[5:0]                ), //i
    .io_axi_b_payload_resp       (io_axi_1_b_payload_resp[1:0]              ), //i
    .io_axi_ar_valid             (txnAgent_1_io_axi_ar_valid                ), //o
    .io_axi_ar_ready             (io_axi_1_ar_ready                         ), //i
    .io_axi_ar_payload_addr      (txnAgent_1_io_axi_ar_payload_addr[63:0]   ), //o
    .io_axi_ar_payload_id        (txnAgent_1_io_axi_ar_payload_id[5:0]      ), //o
    .io_axi_ar_payload_len       (txnAgent_1_io_axi_ar_payload_len[7:0]     ), //o
    .io_axi_ar_payload_size      (txnAgent_1_io_axi_ar_payload_size[2:0]    ), //o
    .io_axi_ar_payload_burst     (txnAgent_1_io_axi_ar_payload_burst[1:0]   ), //o
    .io_axi_r_valid              (io_axi_1_r_valid                          ), //i
    .io_axi_r_ready              (txnAgent_1_io_axi_r_ready                 ), //o
    .io_axi_r_payload_data       (io_axi_1_r_payload_data[511:0]            ), //i
    .io_axi_r_payload_id         (io_axi_1_r_payload_id[5:0]                ), //i
    .io_axi_r_payload_resp       (io_axi_1_r_payload_resp[1:0]              ), //i
    .io_axi_r_payload_last       (io_axi_1_r_payload_last                   ), //i
    .io_ltReq_valid              (txnAgent_1_io_ltReq_valid                 ), //o
    .io_ltReq_ready              (ltMCh_io_lt_1_lkReq_ready                 ), //i
    .io_ltReq_payload_nId        (txnAgent_1_io_ltReq_payload_nId           ), //o
    .io_ltReq_payload_tId        (txnAgent_1_io_ltReq_payload_tId[21:0]     ), //o
    .io_ltReq_payload_tabId      (txnAgent_1_io_ltReq_payload_tabId[2:0]    ), //o
    .io_ltReq_payload_snId       (txnAgent_1_io_ltReq_payload_snId          ), //o
    .io_ltReq_payload_txnId      (txnAgent_1_io_ltReq_payload_txnId[5:0]    ), //o
    .io_ltReq_payload_lkType     (txnAgent_1_io_ltReq_payload_lkType[1:0]   ), //o
    .io_ltReq_payload_lkRelease  (txnAgent_1_io_ltReq_payload_lkRelease     ), //o
    .io_ltReq_payload_txnTimeOut (txnAgent_1_io_ltReq_payload_txnTimeOut    ), //o
    .io_ltReq_payload_txnAbt     (txnAgent_1_io_ltReq_payload_txnAbt        ), //o
    .io_ltReq_payload_lkIdx      (txnAgent_1_io_ltReq_payload_lkIdx[5:0]    ), //o
    .io_ltReq_payload_wLen       (txnAgent_1_io_ltReq_payload_wLen[2:0]     ), //o
    .io_ltResp_valid             (ltMCh_io_lt_1_lkResp_valid                ), //i
    .io_ltResp_ready             (txnAgent_1_io_ltResp_ready                ), //o
    .io_ltResp_payload_nId       (ltMCh_io_lt_1_lkResp_payload_nId          ), //i
    .io_ltResp_payload_tId       (ltMCh_io_lt_1_lkResp_payload_tId[21:0]    ), //i
    .io_ltResp_payload_tabId     (ltMCh_io_lt_1_lkResp_payload_tabId[2:0]   ), //i
    .io_ltResp_payload_snId      (ltMCh_io_lt_1_lkResp_payload_snId         ), //i
    .io_ltResp_payload_txnId     (ltMCh_io_lt_1_lkResp_payload_txnId[5:0]   ), //i
    .io_ltResp_payload_lkType    (ltMCh_io_lt_1_lkResp_payload_lkType[1:0]  ), //i
    .io_ltResp_payload_lkRelease (ltMCh_io_lt_1_lkResp_payload_lkRelease    ), //i
    .io_ltResp_payload_txnAbt    (ltMCh_io_lt_1_lkResp_payload_txnAbt       ), //i
    .io_ltResp_payload_lkIdx     (ltMCh_io_lt_1_lkResp_payload_lkIdx[5:0]   ), //i
    .io_ltResp_payload_wLen      (ltMCh_io_lt_1_lkResp_payload_wLen[2:0]    ), //i
    .io_ltResp_payload_respType  (ltMCh_io_lt_1_lkResp_payload_respType[1:0]), //i
    .io_ltResp_payload_lkWaited  (ltMCh_io_lt_1_lkResp_payload_lkWaited     ), //i
    .clk                         (clk                                       ), //i
    .resetn                      (resetn                                    )  //i
  );
  SendArbiter sendArb (
    .io_lkReqV_0_valid              (txnManAry_0_io_lkReqRmt_valid              ), //i
    .io_lkReqV_0_ready              (sendArb_io_lkReqV_0_ready                  ), //o
    .io_lkReqV_0_payload_nId        (txnManAry_0_io_lkReqRmt_payload_nId        ), //i
    .io_lkReqV_0_payload_tId        (txnManAry_0_io_lkReqRmt_payload_tId[21:0]  ), //i
    .io_lkReqV_0_payload_tabId      (txnManAry_0_io_lkReqRmt_payload_tabId[2:0] ), //i
    .io_lkReqV_0_payload_snId       (txnManAry_0_io_lkReqRmt_payload_snId       ), //i
    .io_lkReqV_0_payload_txnId      (txnManAry_0_io_lkReqRmt_payload_txnId[5:0] ), //i
    .io_lkReqV_0_payload_lkType     (txnManAry_0_io_lkReqRmt_payload_lkType[1:0]), //i
    .io_lkReqV_0_payload_lkRelease  (txnManAry_0_io_lkReqRmt_payload_lkRelease  ), //i
    .io_lkReqV_0_payload_txnTimeOut (txnManAry_0_io_lkReqRmt_payload_txnTimeOut ), //i
    .io_lkReqV_0_payload_txnAbt     (txnManAry_0_io_lkReqRmt_payload_txnAbt     ), //i
    .io_lkReqV_0_payload_lkIdx      (txnManAry_0_io_lkReqRmt_payload_lkIdx[5:0] ), //i
    .io_lkReqV_0_payload_wLen       (txnManAry_0_io_lkReqRmt_payload_wLen[2:0]  ), //i
    .io_wrDataV_0_valid             (txnManAry_0_io_wrRmt_valid                 ), //i
    .io_wrDataV_0_ready             (sendArb_io_wrDataV_0_ready                 ), //o
    .io_wrDataV_0_payload           (txnManAry_0_io_wrRmt_payload[511:0]        ), //i
    .io_sendQ_valid                 (sendArb_io_sendQ_valid                     ), //o
    .io_sendQ_ready                 (io_sendQ_ready                             ), //i
    .io_sendQ_payload               (sendArb_io_sendQ_payload[511:0]            ), //o
    .io_statusVld                   (sendArb_io_statusVld                       ), //o
    .io_nReq                        (sendArb_io_nReq[3:0]                       ), //o
    .io_nWrCmtReq                   (sendArb_io_nWrCmtReq[3:0]                  ), //o
    .io_nRdGetReq                   (sendArb_io_nRdGetReq[3:0]                  ), //o
    .clk                            (clk                                        ), //i
    .resetn                         (resetn                                     )  //i
  );
  RecvDispatcher recvDisp (
    .io_recvQ_valid                 (io_recvQ_valid                             ), //i
    .io_recvQ_ready                 (recvDisp_io_recvQ_ready                    ), //o
    .io_recvQ_payload               (io_recvQ_payload[511:0]                    ), //i
    .io_lkRespV_0_valid             (recvDisp_io_lkRespV_0_valid                ), //o
    .io_lkRespV_0_ready             (txnManAry_0_io_lkRespRmt_ready             ), //i
    .io_lkRespV_0_payload_nId       (recvDisp_io_lkRespV_0_payload_nId          ), //o
    .io_lkRespV_0_payload_tId       (recvDisp_io_lkRespV_0_payload_tId[21:0]    ), //o
    .io_lkRespV_0_payload_tabId     (recvDisp_io_lkRespV_0_payload_tabId[2:0]   ), //o
    .io_lkRespV_0_payload_snId      (recvDisp_io_lkRespV_0_payload_snId         ), //o
    .io_lkRespV_0_payload_txnId     (recvDisp_io_lkRespV_0_payload_txnId[5:0]   ), //o
    .io_lkRespV_0_payload_lkType    (recvDisp_io_lkRespV_0_payload_lkType[1:0]  ), //o
    .io_lkRespV_0_payload_lkRelease (recvDisp_io_lkRespV_0_payload_lkRelease    ), //o
    .io_lkRespV_0_payload_txnAbt    (recvDisp_io_lkRespV_0_payload_txnAbt       ), //o
    .io_lkRespV_0_payload_lkIdx     (recvDisp_io_lkRespV_0_payload_lkIdx[5:0]   ), //o
    .io_lkRespV_0_payload_wLen      (recvDisp_io_lkRespV_0_payload_wLen[2:0]    ), //o
    .io_lkRespV_0_payload_respType  (recvDisp_io_lkRespV_0_payload_respType[1:0]), //o
    .io_lkRespV_0_payload_lkWaited  (recvDisp_io_lkRespV_0_payload_lkWaited     ), //o
    .io_rdDataV_0_valid             (recvDisp_io_rdDataV_0_valid                ), //o
    .io_rdDataV_0_ready             (txnManAry_0_io_rdRmt_ready                 ), //i
    .io_rdDataV_0_payload           (recvDisp_io_rdDataV_0_payload[511:0]       ), //o
    .io_statusVld                   (recvDisp_io_statusVld                      ), //o
    .io_nResp                       (recvDisp_io_nResp[3:0]                     ), //o
    .io_nWrCmtResp                  (recvDisp_io_nWrCmtResp[3:0]                ), //o
    .io_nRdGetResp                  (recvDisp_io_nRdGetResp[3:0]                ), //o
    .clk                            (clk                                        ), //i
    .resetn                         (resetn                                     )  //i
  );
  ReqDispatcher reqDisp (
    .io_reqQ_valid               (io_reqQ_valid                       ), //i
    .io_reqQ_ready               (reqDisp_io_reqQ_ready               ), //o
    .io_reqQ_payload             (io_reqQ_payload[511:0]              ), //i
    .io_lkReq_valid              (reqDisp_io_lkReq_valid              ), //o
    .io_lkReq_ready              (txnAgent_1_io_lkReq_ready           ), //i
    .io_lkReq_payload_nId        (reqDisp_io_lkReq_payload_nId        ), //o
    .io_lkReq_payload_tId        (reqDisp_io_lkReq_payload_tId[21:0]  ), //o
    .io_lkReq_payload_tabId      (reqDisp_io_lkReq_payload_tabId[2:0] ), //o
    .io_lkReq_payload_snId       (reqDisp_io_lkReq_payload_snId       ), //o
    .io_lkReq_payload_txnId      (reqDisp_io_lkReq_payload_txnId[5:0] ), //o
    .io_lkReq_payload_lkType     (reqDisp_io_lkReq_payload_lkType[1:0]), //o
    .io_lkReq_payload_lkRelease  (reqDisp_io_lkReq_payload_lkRelease  ), //o
    .io_lkReq_payload_txnTimeOut (reqDisp_io_lkReq_payload_txnTimeOut ), //o
    .io_lkReq_payload_txnAbt     (reqDisp_io_lkReq_payload_txnAbt     ), //o
    .io_lkReq_payload_lkIdx      (reqDisp_io_lkReq_payload_lkIdx[5:0] ), //o
    .io_lkReq_payload_wLen       (reqDisp_io_lkReq_payload_wLen[2:0]  ), //o
    .io_wrData_valid             (reqDisp_io_wrData_valid             ), //o
    .io_wrData_ready             (txnAgent_1_io_wrData_ready          ), //i
    .io_wrData_payload           (reqDisp_io_wrData_payload[511:0]    ), //o
    .clk                         (clk                                 ), //i
    .resetn                      (resetn                              )  //i
  );
  RespArbiter respArb (
    .io_lkResp_valid             (txnAgent_1_io_lkResp_valid                ), //i
    .io_lkResp_ready             (respArb_io_lkResp_ready                   ), //o
    .io_lkResp_payload_nId       (txnAgent_1_io_lkResp_payload_nId          ), //i
    .io_lkResp_payload_tId       (txnAgent_1_io_lkResp_payload_tId[21:0]    ), //i
    .io_lkResp_payload_tabId     (txnAgent_1_io_lkResp_payload_tabId[2:0]   ), //i
    .io_lkResp_payload_snId      (txnAgent_1_io_lkResp_payload_snId         ), //i
    .io_lkResp_payload_txnId     (txnAgent_1_io_lkResp_payload_txnId[5:0]   ), //i
    .io_lkResp_payload_lkType    (txnAgent_1_io_lkResp_payload_lkType[1:0]  ), //i
    .io_lkResp_payload_lkRelease (txnAgent_1_io_lkResp_payload_lkRelease    ), //i
    .io_lkResp_payload_txnAbt    (txnAgent_1_io_lkResp_payload_txnAbt       ), //i
    .io_lkResp_payload_lkIdx     (txnAgent_1_io_lkResp_payload_lkIdx[5:0]   ), //i
    .io_lkResp_payload_wLen      (txnAgent_1_io_lkResp_payload_wLen[2:0]    ), //i
    .io_lkResp_payload_respType  (txnAgent_1_io_lkResp_payload_respType[1:0]), //i
    .io_lkResp_payload_lkWaited  (txnAgent_1_io_lkResp_payload_lkWaited     ), //i
    .io_rdData_valid             (txnAgent_1_io_rdData_valid                ), //i
    .io_rdData_ready             (respArb_io_rdData_ready                   ), //o
    .io_rdData_payload           (txnAgent_1_io_rdData_payload[511:0]       ), //i
    .io_respQ_valid              (respArb_io_respQ_valid                    ), //o
    .io_respQ_ready              (io_respQ_ready                            ), //i
    .io_respQ_payload            (respArb_io_respQ_payload[511:0]           ), //o
    .clk                         (clk                                       ), //i
    .resetn                      (resetn                                    )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType)
      LkT_rd : txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "insTab";
      default : txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(txnManAry_0_io_lkReqLoc_rData_lkType)
      LkT_rd : txnManAry_0_io_lkReqLoc_rData_lkType_string = "rd    ";
      LkT_wr : txnManAry_0_io_lkReqLoc_rData_lkType_string = "wr    ";
      LkT_raw : txnManAry_0_io_lkReqLoc_rData_lkType_string = "raw   ";
      LkT_insTab : txnManAry_0_io_lkReqLoc_rData_lkType_string = "insTab";
      default : txnManAry_0_io_lkReqLoc_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType)
      LkT_rd : _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType)
      LkT_rd : txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string = "insTab";
      default : txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_rData_lkType)
      LkT_rd : ltMCh_io_lt_0_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltMCh_io_lt_0_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltMCh_io_lt_0_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltMCh_io_lt_0_lkResp_rData_lkType_string = "insTab";
      default : ltMCh_io_lt_0_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_rData_respType)
      LockRespType_grant : ltMCh_io_lt_0_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltMCh_io_lt_0_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltMCh_io_lt_0_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltMCh_io_lt_0_lkResp_rData_respType_string = "release_1";
      default : ltMCh_io_lt_0_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  `endif

  assign io_cmdAxi_0_aw_valid = txnManAry_0_io_cmdAxi_aw_valid;
  assign io_cmdAxi_0_aw_payload_addr = txnManAry_0_io_cmdAxi_aw_payload_addr;
  assign io_cmdAxi_0_aw_payload_id = txnManAry_0_io_cmdAxi_aw_payload_id;
  assign io_cmdAxi_0_aw_payload_len = txnManAry_0_io_cmdAxi_aw_payload_len;
  assign io_cmdAxi_0_aw_payload_size = txnManAry_0_io_cmdAxi_aw_payload_size;
  assign io_cmdAxi_0_aw_payload_burst = txnManAry_0_io_cmdAxi_aw_payload_burst;
  assign io_cmdAxi_0_w_valid = txnManAry_0_io_cmdAxi_w_valid;
  assign io_cmdAxi_0_w_payload_data = txnManAry_0_io_cmdAxi_w_payload_data;
  assign io_cmdAxi_0_w_payload_strb = txnManAry_0_io_cmdAxi_w_payload_strb;
  assign io_cmdAxi_0_w_payload_last = txnManAry_0_io_cmdAxi_w_payload_last;
  assign io_cmdAxi_0_b_ready = txnManAry_0_io_cmdAxi_b_ready;
  assign io_cmdAxi_0_ar_valid = txnManAry_0_io_cmdAxi_ar_valid;
  assign io_cmdAxi_0_ar_payload_addr = txnManAry_0_io_cmdAxi_ar_payload_addr;
  assign io_cmdAxi_0_ar_payload_id = txnManAry_0_io_cmdAxi_ar_payload_id;
  assign io_cmdAxi_0_ar_payload_len = txnManAry_0_io_cmdAxi_ar_payload_len;
  assign io_cmdAxi_0_ar_payload_size = txnManAry_0_io_cmdAxi_ar_payload_size;
  assign io_cmdAxi_0_ar_payload_burst = txnManAry_0_io_cmdAxi_ar_payload_burst;
  assign io_cmdAxi_0_r_ready = txnManAry_0_io_cmdAxi_r_ready;
  assign io_done_0 = txnManAry_0_io_done;
  assign io_cntTxnCmt_0 = txnManAry_0_io_cntTxnCmt;
  assign io_cntTxnAbt_0 = txnManAry_0_io_cntTxnAbt;
  assign io_cntTxnLd_0 = txnManAry_0_io_cntTxnLd;
  assign io_cntClk_0 = txnManAry_0_io_cntClk;
  assign io_cntLockLoc_0 = txnManAry_0_io_cntLockLoc;
  assign io_cntLockRmt_0 = txnManAry_0_io_cntLockRmt;
  assign io_cntLockDenyLoc_0 = txnManAry_0_io_cntLockDenyLoc;
  assign io_cntLockDenyRmt_0 = txnManAry_0_io_cntLockDenyRmt;
  assign io_axi_0_aw_valid = txnManAry_0_io_axi_aw_valid;
  assign io_axi_0_aw_payload_addr = txnManAry_0_io_axi_aw_payload_addr;
  assign io_axi_0_aw_payload_id = txnManAry_0_io_axi_aw_payload_id;
  assign io_axi_0_aw_payload_len = txnManAry_0_io_axi_aw_payload_len;
  assign io_axi_0_aw_payload_size = txnManAry_0_io_axi_aw_payload_size;
  assign io_axi_0_aw_payload_burst = txnManAry_0_io_axi_aw_payload_burst;
  assign io_axi_0_w_valid = txnManAry_0_io_axi_w_valid;
  assign io_axi_0_w_payload_data = txnManAry_0_io_axi_w_payload_data;
  assign io_axi_0_w_payload_strb = txnManAry_0_io_axi_w_payload_strb;
  assign io_axi_0_w_payload_last = txnManAry_0_io_axi_w_payload_last;
  assign io_axi_0_b_ready = txnManAry_0_io_axi_b_ready;
  assign io_axi_0_ar_valid = txnManAry_0_io_axi_ar_valid;
  assign io_axi_0_ar_payload_addr = txnManAry_0_io_axi_ar_payload_addr;
  assign io_axi_0_ar_payload_id = txnManAry_0_io_axi_ar_payload_id;
  assign io_axi_0_ar_payload_len = txnManAry_0_io_axi_ar_payload_len;
  assign io_axi_0_ar_payload_size = txnManAry_0_io_axi_ar_payload_size;
  assign io_axi_0_ar_payload_burst = txnManAry_0_io_axi_ar_payload_burst;
  assign io_axi_0_r_ready = txnManAry_0_io_axi_r_ready;
  assign txnManAry_0_io_lkReqLoc_ready = (! txnManAry_0_io_lkReqLoc_rValid);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_valid = (txnManAry_0_io_lkReqLoc_valid || txnManAry_0_io_lkReqLoc_rValid);
  assign _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_lkType : txnManAry_0_io_lkReqLoc_payload_lkType);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_nId = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_nId : txnManAry_0_io_lkReqLoc_payload_nId);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_tId = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_tId : txnManAry_0_io_lkReqLoc_payload_tId);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_tabId = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_tabId : txnManAry_0_io_lkReqLoc_payload_tabId);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_snId = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_snId : txnManAry_0_io_lkReqLoc_payload_snId);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnId = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_txnId : txnManAry_0_io_lkReqLoc_payload_txnId);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType = _zz_txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkRelease = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_lkRelease : txnManAry_0_io_lkReqLoc_payload_lkRelease);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnTimeOut = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_txnTimeOut : txnManAry_0_io_lkReqLoc_payload_txnTimeOut);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnAbt = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_txnAbt : txnManAry_0_io_lkReqLoc_payload_txnAbt);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkIdx = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_lkIdx : txnManAry_0_io_lkReqLoc_payload_lkIdx);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_payload_wLen = (txnManAry_0_io_lkReqLoc_rValid ? txnManAry_0_io_lkReqLoc_rData_wLen : txnManAry_0_io_lkReqLoc_payload_wLen);
  always @(*) begin
    txnManAry_0_io_lkReqLoc_s2mPipe_ready = txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      txnManAry_0_io_lkReqLoc_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_valid);
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_valid = txnManAry_0_io_lkReqLoc_s2mPipe_rValid;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_nId = txnManAry_0_io_lkReqLoc_s2mPipe_rData_nId;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tId = txnManAry_0_io_lkReqLoc_s2mPipe_rData_tId;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_tabId = txnManAry_0_io_lkReqLoc_s2mPipe_rData_tabId;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_snId = txnManAry_0_io_lkReqLoc_s2mPipe_rData_snId;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnId = txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnId;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkType = txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkRelease = txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkRelease;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnTimeOut = txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnTimeOut;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_txnAbt = txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnAbt;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_lkIdx = txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkIdx;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_payload_wLen = txnManAry_0_io_lkReqLoc_s2mPipe_rData_wLen;
  assign txnManAry_0_io_lkReqLoc_s2mPipe_m2sPipe_ready = ltMCh_io_lt_0_lkReq_ready;
  assign ltMCh_io_lt_0_lkResp_ready = (! ltMCh_io_lt_0_lkResp_rValid);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_valid = (ltMCh_io_lt_0_lkResp_valid || ltMCh_io_lt_0_lkResp_rValid);
  assign _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_lkType : ltMCh_io_lt_0_lkResp_payload_lkType);
  assign _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_respType : ltMCh_io_lt_0_lkResp_payload_respType);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_nId = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_nId : ltMCh_io_lt_0_lkResp_payload_nId);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_tId = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_tId : ltMCh_io_lt_0_lkResp_payload_tId);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_tabId = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_tabId : ltMCh_io_lt_0_lkResp_payload_tabId);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_snId = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_snId : ltMCh_io_lt_0_lkResp_payload_snId);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnId = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_txnId : ltMCh_io_lt_0_lkResp_payload_txnId);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType = _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkRelease = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_lkRelease : ltMCh_io_lt_0_lkResp_payload_lkRelease);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnAbt = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_txnAbt : ltMCh_io_lt_0_lkResp_payload_txnAbt);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkIdx = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_lkIdx : ltMCh_io_lt_0_lkResp_payload_lkIdx);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_wLen = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_wLen : ltMCh_io_lt_0_lkResp_payload_wLen);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType = _zz_ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkWaited = (ltMCh_io_lt_0_lkResp_rValid ? ltMCh_io_lt_0_lkResp_rData_lkWaited : ltMCh_io_lt_0_lkResp_payload_lkWaited);
  always @(*) begin
    ltMCh_io_lt_0_lkResp_s2mPipe_ready = ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      ltMCh_io_lt_0_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_valid);
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_valid = ltMCh_io_lt_0_lkResp_s2mPipe_rValid;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_nId = ltMCh_io_lt_0_lkResp_s2mPipe_rData_nId;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tId = ltMCh_io_lt_0_lkResp_s2mPipe_rData_tId;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_tabId = ltMCh_io_lt_0_lkResp_s2mPipe_rData_tabId;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_snId = ltMCh_io_lt_0_lkResp_s2mPipe_rData_snId;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnId = ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnId;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkType = ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkRelease;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnAbt;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkIdx;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_wLen = ltMCh_io_lt_0_lkResp_s2mPipe_rData_wLen;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_respType = ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkWaited;
  assign ltMCh_io_lt_0_lkResp_s2mPipe_m2sPipe_ready = txnManAry_0_io_lkRespLoc_ready;
  assign io_sendQ_valid = sendArb_io_sendQ_valid;
  assign io_sendQ_payload = sendArb_io_sendQ_payload;
  assign io_recvQ_ready = recvDisp_io_recvQ_ready;
  assign io_reqQ_ready = reqDisp_io_reqQ_ready;
  assign io_respQ_valid = respArb_io_respQ_valid;
  assign io_respQ_payload = respArb_io_respQ_payload;
  assign io_sendStatusVld = sendArb_io_statusVld;
  assign io_nReq = sendArb_io_nReq;
  assign io_nWrCmtReq = sendArb_io_nWrCmtReq;
  assign io_nRdGetReq = sendArb_io_nRdGetReq;
  assign io_recvStatusVld = recvDisp_io_statusVld;
  assign io_nResp = recvDisp_io_nResp;
  assign io_nWrCmtResp = recvDisp_io_nWrCmtResp;
  assign io_nRdGetResp = recvDisp_io_nRdGetResp;
  assign io_axi_1_aw_valid = txnAgent_1_io_axi_aw_valid;
  assign io_axi_1_aw_payload_addr = txnAgent_1_io_axi_aw_payload_addr;
  assign io_axi_1_aw_payload_id = txnAgent_1_io_axi_aw_payload_id;
  assign io_axi_1_aw_payload_len = txnAgent_1_io_axi_aw_payload_len;
  assign io_axi_1_aw_payload_size = txnAgent_1_io_axi_aw_payload_size;
  assign io_axi_1_aw_payload_burst = txnAgent_1_io_axi_aw_payload_burst;
  assign io_axi_1_w_valid = txnAgent_1_io_axi_w_valid;
  assign io_axi_1_w_payload_data = txnAgent_1_io_axi_w_payload_data;
  assign io_axi_1_w_payload_strb = txnAgent_1_io_axi_w_payload_strb;
  assign io_axi_1_w_payload_last = txnAgent_1_io_axi_w_payload_last;
  assign io_axi_1_b_ready = txnAgent_1_io_axi_b_ready;
  assign io_axi_1_ar_valid = txnAgent_1_io_axi_ar_valid;
  assign io_axi_1_ar_payload_addr = txnAgent_1_io_axi_ar_payload_addr;
  assign io_axi_1_ar_payload_id = txnAgent_1_io_axi_ar_payload_id;
  assign io_axi_1_ar_payload_len = txnAgent_1_io_axi_ar_payload_len;
  assign io_axi_1_ar_payload_size = txnAgent_1_io_axi_ar_payload_size;
  assign io_axi_1_ar_payload_burst = txnAgent_1_io_axi_ar_payload_burst;
  assign io_axi_1_r_ready = txnAgent_1_io_axi_r_ready;
  always @(posedge clk) begin
    if(!resetn) begin
      txnManAry_0_io_lkReqLoc_rValid <= 1'b0;
      txnManAry_0_io_lkReqLoc_s2mPipe_rValid <= 1'b0;
      ltMCh_io_lt_0_lkResp_rValid <= 1'b0;
      ltMCh_io_lt_0_lkResp_s2mPipe_rValid <= 1'b0;
    end else begin
      if(txnManAry_0_io_lkReqLoc_valid) begin
        txnManAry_0_io_lkReqLoc_rValid <= 1'b1;
      end
      if(txnManAry_0_io_lkReqLoc_s2mPipe_ready) begin
        txnManAry_0_io_lkReqLoc_rValid <= 1'b0;
      end
      if(txnManAry_0_io_lkReqLoc_s2mPipe_ready) begin
        txnManAry_0_io_lkReqLoc_s2mPipe_rValid <= txnManAry_0_io_lkReqLoc_s2mPipe_valid;
      end
      if(ltMCh_io_lt_0_lkResp_valid) begin
        ltMCh_io_lt_0_lkResp_rValid <= 1'b1;
      end
      if(ltMCh_io_lt_0_lkResp_s2mPipe_ready) begin
        ltMCh_io_lt_0_lkResp_rValid <= 1'b0;
      end
      if(ltMCh_io_lt_0_lkResp_s2mPipe_ready) begin
        ltMCh_io_lt_0_lkResp_s2mPipe_rValid <= ltMCh_io_lt_0_lkResp_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(txnManAry_0_io_lkReqLoc_ready) begin
      txnManAry_0_io_lkReqLoc_rData_nId <= txnManAry_0_io_lkReqLoc_payload_nId;
      txnManAry_0_io_lkReqLoc_rData_tId <= txnManAry_0_io_lkReqLoc_payload_tId;
      txnManAry_0_io_lkReqLoc_rData_tabId <= txnManAry_0_io_lkReqLoc_payload_tabId;
      txnManAry_0_io_lkReqLoc_rData_snId <= txnManAry_0_io_lkReqLoc_payload_snId;
      txnManAry_0_io_lkReqLoc_rData_txnId <= txnManAry_0_io_lkReqLoc_payload_txnId;
      txnManAry_0_io_lkReqLoc_rData_lkType <= txnManAry_0_io_lkReqLoc_payload_lkType;
      txnManAry_0_io_lkReqLoc_rData_lkRelease <= txnManAry_0_io_lkReqLoc_payload_lkRelease;
      txnManAry_0_io_lkReqLoc_rData_txnTimeOut <= txnManAry_0_io_lkReqLoc_payload_txnTimeOut;
      txnManAry_0_io_lkReqLoc_rData_txnAbt <= txnManAry_0_io_lkReqLoc_payload_txnAbt;
      txnManAry_0_io_lkReqLoc_rData_lkIdx <= txnManAry_0_io_lkReqLoc_payload_lkIdx;
      txnManAry_0_io_lkReqLoc_rData_wLen <= txnManAry_0_io_lkReqLoc_payload_wLen;
    end
    if(txnManAry_0_io_lkReqLoc_s2mPipe_ready) begin
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_nId <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_nId;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_tId <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_tId;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_tabId <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_tabId;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_snId <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_snId;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnId <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnId;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkType <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkType;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkRelease <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkRelease;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnTimeOut <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnTimeOut;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_txnAbt <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_txnAbt;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_lkIdx <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_lkIdx;
      txnManAry_0_io_lkReqLoc_s2mPipe_rData_wLen <= txnManAry_0_io_lkReqLoc_s2mPipe_payload_wLen;
    end
    if(ltMCh_io_lt_0_lkResp_ready) begin
      ltMCh_io_lt_0_lkResp_rData_nId <= ltMCh_io_lt_0_lkResp_payload_nId;
      ltMCh_io_lt_0_lkResp_rData_tId <= ltMCh_io_lt_0_lkResp_payload_tId;
      ltMCh_io_lt_0_lkResp_rData_tabId <= ltMCh_io_lt_0_lkResp_payload_tabId;
      ltMCh_io_lt_0_lkResp_rData_snId <= ltMCh_io_lt_0_lkResp_payload_snId;
      ltMCh_io_lt_0_lkResp_rData_txnId <= ltMCh_io_lt_0_lkResp_payload_txnId;
      ltMCh_io_lt_0_lkResp_rData_lkType <= ltMCh_io_lt_0_lkResp_payload_lkType;
      ltMCh_io_lt_0_lkResp_rData_lkRelease <= ltMCh_io_lt_0_lkResp_payload_lkRelease;
      ltMCh_io_lt_0_lkResp_rData_txnAbt <= ltMCh_io_lt_0_lkResp_payload_txnAbt;
      ltMCh_io_lt_0_lkResp_rData_lkIdx <= ltMCh_io_lt_0_lkResp_payload_lkIdx;
      ltMCh_io_lt_0_lkResp_rData_wLen <= ltMCh_io_lt_0_lkResp_payload_wLen;
      ltMCh_io_lt_0_lkResp_rData_respType <= ltMCh_io_lt_0_lkResp_payload_respType;
      ltMCh_io_lt_0_lkResp_rData_lkWaited <= ltMCh_io_lt_0_lkResp_payload_lkWaited;
    end
    if(ltMCh_io_lt_0_lkResp_s2mPipe_ready) begin
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_nId <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_nId;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_tId <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_tId;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_tabId <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_tabId;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_snId <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_snId;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnId <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnId;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkType <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkType;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkRelease <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkRelease;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_txnAbt <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_txnAbt;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkIdx <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkIdx;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_wLen <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_wLen;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_respType <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_respType;
      ltMCh_io_lt_0_lkResp_s2mPipe_rData_lkWaited <= ltMCh_io_lt_0_lkResp_s2mPipe_payload_lkWaited;
    end
  end


endmodule

module StreamDemux_6 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [42:0]   io_input_payload_data,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [42:0]   io_outputs_0_payload_data,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [42:0]   io_outputs_1_payload_data
);

  wire                when_Stream_l881;
  wire                when_Stream_l881_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l881) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l881_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_data = io_input_payload_data;
  assign when_Stream_l881 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l881) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_data = io_input_payload_data;
  assign when_Stream_l881_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l881_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module StreamDemux_5 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [511:0]  io_input_payload_tdata,
  input      [63:0]   io_input_payload_tkeep,
  input               io_input_payload_tlast,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [511:0]  io_outputs_0_payload_tdata,
  output     [63:0]   io_outputs_0_payload_tkeep,
  output              io_outputs_0_payload_tlast,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [511:0]  io_outputs_1_payload_tdata,
  output     [63:0]   io_outputs_1_payload_tkeep,
  output              io_outputs_1_payload_tlast
);

  wire                when_Stream_l881;
  wire                when_Stream_l881_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l881) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l881_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_tdata = io_input_payload_tdata;
  assign io_outputs_0_payload_tkeep = io_input_payload_tkeep;
  assign io_outputs_0_payload_tlast = io_input_payload_tlast;
  assign when_Stream_l881 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l881) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_tdata = io_input_payload_tdata;
  assign io_outputs_1_payload_tkeep = io_input_payload_tkeep;
  assign io_outputs_1_payload_tlast = io_input_payload_tlast;
  assign when_Stream_l881_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l881_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

//StreamDemux_3 replaced by StreamDemux_3

//StreamFifo_7 replaced by StreamFifo_7

module StreamMux_1 (
  input      [0:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [511:0]  io_inputs_0_payload_tdata,
  input      [63:0]   io_inputs_0_payload_tkeep,
  input               io_inputs_0_payload_tlast,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [511:0]  io_inputs_1_payload_tdata,
  input      [63:0]   io_inputs_1_payload_tkeep,
  input               io_inputs_1_payload_tlast,
  output              io_output_valid,
  input               io_output_ready,
  output     [511:0]  io_output_payload_tdata,
  output     [63:0]   io_output_payload_tkeep,
  output              io_output_payload_tlast
);

  reg                 _zz_io_output_valid;
  reg        [511:0]  _zz_io_output_payload_tdata;
  reg        [63:0]   _zz_io_output_payload_tkeep;
  reg                 _zz_io_output_payload_tlast;

  always @(*) begin
    case(io_select)
      1'b0 : begin
        _zz_io_output_valid = io_inputs_0_valid;
        _zz_io_output_payload_tdata = io_inputs_0_payload_tdata;
        _zz_io_output_payload_tkeep = io_inputs_0_payload_tkeep;
        _zz_io_output_payload_tlast = io_inputs_0_payload_tlast;
      end
      default : begin
        _zz_io_output_valid = io_inputs_1_valid;
        _zz_io_output_payload_tdata = io_inputs_1_payload_tdata;
        _zz_io_output_payload_tkeep = io_inputs_1_payload_tkeep;
        _zz_io_output_payload_tlast = io_inputs_1_payload_tlast;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 1'b0) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 1'b1) && io_output_ready);
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_tdata = _zz_io_output_payload_tdata;
  assign io_output_payload_tkeep = _zz_io_output_payload_tkeep;
  assign io_output_payload_tlast = _zz_io_output_payload_tlast;

endmodule

module StreamDemux_3 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [95:0]   io_input_payload_data,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [95:0]   io_outputs_0_payload_data,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [95:0]   io_outputs_1_payload_data
);

  wire                when_Stream_l881;
  wire                when_Stream_l881_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l881) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l881_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_data = io_input_payload_data;
  assign when_Stream_l881 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l881) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_data = io_input_payload_data;
  assign when_Stream_l881_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l881_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module StreamMux (
  input      [0:0]    io_select,
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [543:0]  io_inputs_0_payload_data,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [543:0]  io_inputs_1_payload_data,
  output              io_output_valid,
  input               io_output_ready,
  output     [543:0]  io_output_payload_data
);

  reg                 _zz_io_output_valid;
  reg        [543:0]  _zz_io_output_payload_data;

  always @(*) begin
    case(io_select)
      1'b0 : begin
        _zz_io_output_valid = io_inputs_0_valid;
        _zz_io_output_payload_data = io_inputs_0_payload_data;
      end
      default : begin
        _zz_io_output_valid = io_inputs_1_valid;
        _zz_io_output_payload_data = io_inputs_1_payload_data;
      end
    endcase
  end

  assign io_inputs_0_ready = ((io_select == 1'b0) && io_output_ready);
  assign io_inputs_1_ready = ((io_select == 1'b1) && io_output_ready);
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_data = _zz_io_output_payload_data;

endmodule

//StreamFifo_7 replaced by StreamFifo_7

module StreamFifo_7 (
  input               io_push_valid,
  output              io_push_ready,
  input      [0:0]    io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [0:0]    io_pop_payload,
  input               io_flush,
  output     [5:0]    io_occupancy,
  output     [5:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [0:0]    _zz_logic_ram_port0;
  wire       [4:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [4:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [0:0]    _zz_logic_ram_port_1;
  wire       [4:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [4:0]    logic_pushPtr_valueNext;
  reg        [4:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [4:0]    logic_popPtr_valueNext;
  reg        [4:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1075;
  wire       [4:0]    logic_ptrDif;
  reg [0:0] logic_ram [0:31];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {4'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {4'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  assign _zz_logic_ram_port_1 = io_push_payload;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 5'h1f);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 5'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 5'h1f);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 5'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 5'h0;
      logic_popPtr_value <= 5'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1075) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

//StreamFifo_3 replaced by StreamFifo_3

//StreamFifo_3 replaced by StreamFifo_3

//StreamFifo_3 replaced by StreamFifo_3

module StreamFifo_3 (
  input               io_push_valid,
  output              io_push_ready,
  input      [511:0]  io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [511:0]  io_pop_payload,
  input               io_flush,
  output     [9:0]    io_occupancy,
  output     [9:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [511:0]  _zz_logic_ram_port0;
  wire       [8:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [8:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [8:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [8:0]    logic_pushPtr_valueNext;
  reg        [8:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [8:0]    logic_popPtr_valueNext;
  reg        [8:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1075;
  wire       [8:0]    logic_ptrDif;
  reg [511:0] logic_ram [0:511];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {8'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {8'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 9'h1ff);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 9'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 9'h1ff);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 9'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 9'h0;
      logic_popPtr_value <= 9'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1075) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module RespArbiter (
  input               io_lkResp_valid,
  output reg          io_lkResp_ready,
  input      [0:0]    io_lkResp_payload_nId,
  input      [21:0]   io_lkResp_payload_tId,
  input      [2:0]    io_lkResp_payload_tabId,
  input      [0:0]    io_lkResp_payload_snId,
  input      [5:0]    io_lkResp_payload_txnId,
  input      [1:0]    io_lkResp_payload_lkType,
  input               io_lkResp_payload_lkRelease,
  input               io_lkResp_payload_txnAbt,
  input      [5:0]    io_lkResp_payload_lkIdx,
  input      [2:0]    io_lkResp_payload_wLen,
  input      [1:0]    io_lkResp_payload_respType,
  input               io_lkResp_payload_lkWaited,
  input               io_rdData_valid,
  output reg          io_rdData_ready,
  input      [511:0]  io_rdData_payload,
  output reg          io_respQ_valid,
  input               io_respQ_ready,
  output reg [511:0]  io_respQ_payload,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam fsm_enumDef_4_BOOT = 2'd0;
  localparam fsm_enumDef_4_LKRESP = 2'd1;
  localparam fsm_enumDef_4_RDDATA = 2'd2;

  wire                _zz_when;
  wire       [48:0]   _zz_io_respQ_payload;
  wire       [21:0]   _zz_io_respQ_payload_1;
  wire       [0:0]    _zz_io_respQ_payload_2;
  wire       [11:0]   _zz_cntBeat;
  wire       [7:0]    _zz_cntBeat_1;
  reg        [11:0]   cntBeat;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 io_lkResp_slowdown_x1_valid;
  wire                io_lkResp_slowdown_x1_ready;
  wire       [0:0]    io_lkResp_slowdown_x1_payload_0_nId;
  wire       [21:0]   io_lkResp_slowdown_x1_payload_0_tId;
  wire       [2:0]    io_lkResp_slowdown_x1_payload_0_tabId;
  wire       [0:0]    io_lkResp_slowdown_x1_payload_0_snId;
  wire       [5:0]    io_lkResp_slowdown_x1_payload_0_txnId;
  wire       [1:0]    io_lkResp_slowdown_x1_payload_0_lkType;
  wire                io_lkResp_slowdown_x1_payload_0_lkRelease;
  wire                io_lkResp_slowdown_x1_payload_0_txnAbt;
  wire       [5:0]    io_lkResp_slowdown_x1_payload_0_lkIdx;
  wire       [2:0]    io_lkResp_slowdown_x1_payload_0_wLen;
  wire       [1:0]    io_lkResp_slowdown_x1_payload_0_respType;
  wire                io_lkResp_slowdown_x1_payload_0_lkWaited;
  wire                io_lkResp_fire;
  wire                _zz_io_lkResp_slowdown_x1_ready;
  wire                fsm_lkRespSlowDown_valid;
  wire                fsm_lkRespSlowDown_ready;
  wire       [0:0]    fsm_lkRespSlowDown_payload_0_nId;
  wire       [21:0]   fsm_lkRespSlowDown_payload_0_tId;
  wire       [2:0]    fsm_lkRespSlowDown_payload_0_tabId;
  wire       [0:0]    fsm_lkRespSlowDown_payload_0_snId;
  wire       [5:0]    fsm_lkRespSlowDown_payload_0_txnId;
  wire       [1:0]    fsm_lkRespSlowDown_payload_0_lkType;
  wire                fsm_lkRespSlowDown_payload_0_lkRelease;
  wire                fsm_lkRespSlowDown_payload_0_txnAbt;
  wire       [5:0]    fsm_lkRespSlowDown_payload_0_lkIdx;
  wire       [2:0]    fsm_lkRespSlowDown_payload_0_wLen;
  wire       [1:0]    fsm_lkRespSlowDown_payload_0_respType;
  wire                fsm_lkRespSlowDown_payload_0_lkWaited;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                _zz_when_NetArb_l300;
  wire                io_lkResp_fire_1;
  wire                when_NetArb_l300;
  wire                io_respQ_fire;
  wire                when_NetArb_l306;
  wire                io_respQ_fire_1;
  wire                when_NetArb_l316;
  `ifndef SYNTHESIS
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] io_lkResp_slowdown_x1_payload_0_lkType_string;
  reg [71:0] io_lkResp_slowdown_x1_payload_0_respType_string;
  reg [47:0] fsm_lkRespSlowDown_payload_0_lkType_string;
  reg [71:0] fsm_lkRespSlowDown_payload_0_respType_string;
  reg [47:0] fsm_stateReg_string;
  reg [47:0] fsm_stateNext_string;
  `endif


  assign _zz_when = 1'b1;
  assign _zz_io_respQ_payload = {fsm_lkRespSlowDown_payload_0_lkWaited,{fsm_lkRespSlowDown_payload_0_respType,{fsm_lkRespSlowDown_payload_0_wLen,{fsm_lkRespSlowDown_payload_0_lkIdx,{fsm_lkRespSlowDown_payload_0_txnAbt,{fsm_lkRespSlowDown_payload_0_lkRelease,{fsm_lkRespSlowDown_payload_0_lkType,{fsm_lkRespSlowDown_payload_0_txnId,{fsm_lkRespSlowDown_payload_0_snId,{fsm_lkRespSlowDown_payload_0_tabId,{_zz_io_respQ_payload_1,_zz_io_respQ_payload_2}}}}}}}}}}};
  assign _zz_cntBeat_1 = ({7'd0,1'b1} <<< io_lkResp_payload_wLen);
  assign _zz_cntBeat = {4'd0, _zz_cntBeat_1};
  assign _zz_io_respQ_payload_1 = fsm_lkRespSlowDown_payload_0_tId;
  assign _zz_io_respQ_payload_2 = fsm_lkRespSlowDown_payload_0_nId;
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_slowdown_x1_payload_0_lkType)
      LkT_rd : io_lkResp_slowdown_x1_payload_0_lkType_string = "rd    ";
      LkT_wr : io_lkResp_slowdown_x1_payload_0_lkType_string = "wr    ";
      LkT_raw : io_lkResp_slowdown_x1_payload_0_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_slowdown_x1_payload_0_lkType_string = "insTab";
      default : io_lkResp_slowdown_x1_payload_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_slowdown_x1_payload_0_respType)
      LockRespType_grant : io_lkResp_slowdown_x1_payload_0_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_slowdown_x1_payload_0_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_slowdown_x1_payload_0_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_slowdown_x1_payload_0_respType_string = "release_1";
      default : io_lkResp_slowdown_x1_payload_0_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_lkRespSlowDown_payload_0_lkType)
      LkT_rd : fsm_lkRespSlowDown_payload_0_lkType_string = "rd    ";
      LkT_wr : fsm_lkRespSlowDown_payload_0_lkType_string = "wr    ";
      LkT_raw : fsm_lkRespSlowDown_payload_0_lkType_string = "raw   ";
      LkT_insTab : fsm_lkRespSlowDown_payload_0_lkType_string = "insTab";
      default : fsm_lkRespSlowDown_payload_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_lkRespSlowDown_payload_0_respType)
      LockRespType_grant : fsm_lkRespSlowDown_payload_0_respType_string = "grant    ";
      LockRespType_abort : fsm_lkRespSlowDown_payload_0_respType_string = "abort    ";
      LockRespType_waiting : fsm_lkRespSlowDown_payload_0_respType_string = "waiting  ";
      LockRespType_release_1 : fsm_lkRespSlowDown_payload_0_respType_string = "release_1";
      default : fsm_lkRespSlowDown_payload_0_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_4_BOOT : fsm_stateReg_string = "BOOT  ";
      fsm_enumDef_4_LKRESP : fsm_stateReg_string = "LKRESP";
      fsm_enumDef_4_RDDATA : fsm_stateReg_string = "RDDATA";
      default : fsm_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_4_BOOT : fsm_stateNext_string = "BOOT  ";
      fsm_enumDef_4_LKRESP : fsm_stateNext_string = "LKRESP";
      fsm_enumDef_4_RDDATA : fsm_stateNext_string = "RDDATA";
      default : fsm_stateNext_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_rdData_ready = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_4_LKRESP : begin
      end
      fsm_enumDef_4_RDDATA : begin
        io_rdData_ready = io_respQ_ready;
      end
      default : begin
      end
    endcase
  end

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_4_LKRESP : begin
      end
      fsm_enumDef_4_RDDATA : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  assign io_lkResp_slowdown_x1_payload_0_nId = io_lkResp_payload_nId;
  assign io_lkResp_slowdown_x1_payload_0_tId = io_lkResp_payload_tId;
  assign io_lkResp_slowdown_x1_payload_0_tabId = io_lkResp_payload_tabId;
  assign io_lkResp_slowdown_x1_payload_0_snId = io_lkResp_payload_snId;
  assign io_lkResp_slowdown_x1_payload_0_txnId = io_lkResp_payload_txnId;
  assign io_lkResp_slowdown_x1_payload_0_lkType = io_lkResp_payload_lkType;
  assign io_lkResp_slowdown_x1_payload_0_lkRelease = io_lkResp_payload_lkRelease;
  assign io_lkResp_slowdown_x1_payload_0_txnAbt = io_lkResp_payload_txnAbt;
  assign io_lkResp_slowdown_x1_payload_0_lkIdx = io_lkResp_payload_lkIdx;
  assign io_lkResp_slowdown_x1_payload_0_wLen = io_lkResp_payload_wLen;
  assign io_lkResp_slowdown_x1_payload_0_respType = io_lkResp_payload_respType;
  assign io_lkResp_slowdown_x1_payload_0_lkWaited = io_lkResp_payload_lkWaited;
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  always @(*) begin
    if(_zz_when) begin
      io_lkResp_ready = io_lkResp_slowdown_x1_ready;
    end else begin
      io_lkResp_ready = 1'b1;
    end
  end

  always @(*) begin
    if(_zz_when) begin
      io_lkResp_slowdown_x1_valid = io_lkResp_valid;
    end else begin
      io_lkResp_slowdown_x1_valid = 1'b0;
    end
  end

  assign fsm_lkRespSlowDown_valid = (io_lkResp_slowdown_x1_valid && _zz_io_lkResp_slowdown_x1_ready);
  assign io_lkResp_slowdown_x1_ready = (fsm_lkRespSlowDown_ready && _zz_io_lkResp_slowdown_x1_ready);
  assign fsm_lkRespSlowDown_payload_0_nId = io_lkResp_slowdown_x1_payload_0_nId;
  assign fsm_lkRespSlowDown_payload_0_tId = io_lkResp_slowdown_x1_payload_0_tId;
  assign fsm_lkRespSlowDown_payload_0_tabId = io_lkResp_slowdown_x1_payload_0_tabId;
  assign fsm_lkRespSlowDown_payload_0_snId = io_lkResp_slowdown_x1_payload_0_snId;
  assign fsm_lkRespSlowDown_payload_0_txnId = io_lkResp_slowdown_x1_payload_0_txnId;
  assign fsm_lkRespSlowDown_payload_0_lkType = io_lkResp_slowdown_x1_payload_0_lkType;
  assign fsm_lkRespSlowDown_payload_0_lkRelease = io_lkResp_slowdown_x1_payload_0_lkRelease;
  assign fsm_lkRespSlowDown_payload_0_txnAbt = io_lkResp_slowdown_x1_payload_0_txnAbt;
  assign fsm_lkRespSlowDown_payload_0_lkIdx = io_lkResp_slowdown_x1_payload_0_lkIdx;
  assign fsm_lkRespSlowDown_payload_0_wLen = io_lkResp_slowdown_x1_payload_0_wLen;
  assign fsm_lkRespSlowDown_payload_0_respType = io_lkResp_slowdown_x1_payload_0_respType;
  assign fsm_lkRespSlowDown_payload_0_lkWaited = io_lkResp_slowdown_x1_payload_0_lkWaited;
  always @(*) begin
    io_respQ_valid = fsm_lkRespSlowDown_valid;
    case(fsm_stateReg)
      fsm_enumDef_4_LKRESP : begin
      end
      fsm_enumDef_4_RDDATA : begin
        io_respQ_valid = io_rdData_valid;
      end
      default : begin
      end
    endcase
  end

  assign fsm_lkRespSlowDown_ready = io_respQ_ready;
  always @(*) begin
    io_respQ_payload = {463'd0, _zz_io_respQ_payload};
    case(fsm_stateReg)
      fsm_enumDef_4_LKRESP : begin
      end
      fsm_enumDef_4_RDDATA : begin
        io_respQ_payload = io_rdData_payload;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_4_LKRESP : begin
        if(io_respQ_fire) begin
          if(when_NetArb_l306) begin
            fsm_stateNext = fsm_enumDef_4_RDDATA;
          end
        end
      end
      fsm_enumDef_4_RDDATA : begin
        if(io_respQ_fire_1) begin
          if(when_NetArb_l316) begin
            fsm_stateNext = fsm_enumDef_4_LKRESP;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_4_LKRESP;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_4_BOOT;
    end
  end

  assign _zz_when_NetArb_l300 = (((! io_lkResp_payload_lkRelease) && ((io_lkResp_payload_lkType == LkT_rd) || (io_lkResp_payload_lkType == LkT_raw))) && (io_lkResp_payload_respType == LockRespType_grant));
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign when_NetArb_l300 = (io_lkResp_fire_1 && _zz_when_NetArb_l300);
  assign io_respQ_fire = (io_respQ_valid && io_respQ_ready);
  assign when_NetArb_l306 = ((cntBeat != 12'h0) || _zz_when_NetArb_l300);
  assign io_respQ_fire_1 = (io_respQ_valid && io_respQ_ready);
  assign when_NetArb_l316 = (cntBeat == 12'h001);
  assign _zz_io_lkResp_slowdown_x1_ready = (fsm_stateReg == fsm_enumDef_4_LKRESP);
  always @(posedge clk) begin
    if(!resetn) begin
      cntBeat <= 12'h0;
      fsm_stateReg <= fsm_enumDef_4_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_4_LKRESP : begin
          if(when_NetArb_l300) begin
            cntBeat <= (cntBeat + _zz_cntBeat);
          end
        end
        fsm_enumDef_4_RDDATA : begin
          if(io_respQ_fire_1) begin
            cntBeat <= (cntBeat - 12'h001);
            if(when_NetArb_l316) begin
              cntBeat <= 12'h0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end


endmodule

module ReqDispatcher (
  input               io_reqQ_valid,
  output reg          io_reqQ_ready,
  input      [511:0]  io_reqQ_payload,
  output reg          io_lkReq_valid,
  input               io_lkReq_ready,
  output     [0:0]    io_lkReq_payload_nId,
  output     [21:0]   io_lkReq_payload_tId,
  output     [2:0]    io_lkReq_payload_tabId,
  output     [0:0]    io_lkReq_payload_snId,
  output     [5:0]    io_lkReq_payload_txnId,
  output     [1:0]    io_lkReq_payload_lkType,
  output              io_lkReq_payload_lkRelease,
  output              io_lkReq_payload_txnTimeOut,
  output              io_lkReq_payload_txnAbt,
  output     [5:0]    io_lkReq_payload_lkIdx,
  output     [2:0]    io_lkReq_payload_wLen,
  output reg          io_wrData_valid,
  input               io_wrData_ready,
  output reg [511:0]  io_wrData_payload,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam fsm_enumDef_3_BOOT = 2'd0;
  localparam fsm_enumDef_3_LKREQ = 2'd1;
  localparam fsm_enumDef_3_LKREQFIRE = 2'd2;
  localparam fsm_enumDef_3_WRDATA = 2'd3;

  wire       [46:0]   _zz_fsm_lkReqBitV_0;
  wire       [0:0]    _zz_fsm_rMskWr_ohFirst_masked;
  wire       [7:0]    _zz_when_NetArb_l261;
  wire       [7:0]    _zz_when_NetArb_l261_1;
  reg        [7:0]    cntBeat;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 fsm_cntFire_willIncrement;
  wire                fsm_cntFire_willClear;
  wire                fsm_cntFire_willOverflowIfInc;
  wire                fsm_cntFire_willOverflow;
  reg        [0:0]    fsm_rLkReq_0_nId;
  reg        [21:0]   fsm_rLkReq_0_tId;
  reg        [2:0]    fsm_rLkReq_0_tabId;
  reg        [0:0]    fsm_rLkReq_0_snId;
  reg        [5:0]    fsm_rLkReq_0_txnId;
  reg        [1:0]    fsm_rLkReq_0_lkType;
  reg                 fsm_rLkReq_0_lkRelease;
  reg                 fsm_rLkReq_0_txnTimeOut;
  reg                 fsm_rLkReq_0_txnAbt;
  reg        [5:0]    fsm_rLkReq_0_lkIdx;
  reg        [2:0]    fsm_rLkReq_0_wLen;
  wire       [46:0]   fsm_lkReqBitV_0;
  wire       [0:0]    fsm_lkReqV_0_nId;
  wire       [21:0]   fsm_lkReqV_0_tId;
  wire       [2:0]    fsm_lkReqV_0_tabId;
  wire       [0:0]    fsm_lkReqV_0_snId;
  wire       [5:0]    fsm_lkReqV_0_txnId;
  wire       [1:0]    fsm_lkReqV_0_lkType;
  wire                fsm_lkReqV_0_lkRelease;
  wire                fsm_lkReqV_0_txnTimeOut;
  wire                fsm_lkReqV_0_txnAbt;
  wire       [5:0]    fsm_lkReqV_0_lkIdx;
  wire       [2:0]    fsm_lkReqV_0_wLen;
  wire       [1:0]    _zz_fsm_lkReqV_0_lkType;
  reg        [0:0]    fsm_rMskWr;
  wire       [0:0]    fsm_MskWr;
  wire       [1:0]    _zz_io_lkReq_payload_lkType;
  wire                _zz_io_reqQ_ready;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                io_reqQ_fire;
  wire                io_lkReq_fire;
  wire                switch_NetArb_l241;
  wire       [0:0]    fsm_rMskWr_ohFirst_input;
  wire       [0:0]    fsm_rMskWr_ohFirst_masked;
  wire       [0:0]    fsm_rMskWr_ohFirst_value;
  reg        [0:0]    _zz_when_NetArb_l265;
  wire                io_reqQ_fire_1;
  wire                when_NetArb_l261;
  wire                when_NetArb_l265;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] fsm_rLkReq_0_lkType_string;
  reg [47:0] fsm_lkReqV_0_lkType_string;
  reg [47:0] _zz_fsm_lkReqV_0_lkType_string;
  reg [47:0] _zz_io_lkReq_payload_lkType_string;
  reg [71:0] fsm_stateReg_string;
  reg [71:0] fsm_stateNext_string;
  `endif


  assign _zz_fsm_lkReqBitV_0 = io_reqQ_payload[46 : 0];
  assign _zz_fsm_rMskWr_ohFirst_masked = (fsm_rMskWr_ohFirst_input - 1'b1);
  assign _zz_when_NetArb_l261 = (_zz_when_NetArb_l261_1 - 8'h01);
  assign _zz_when_NetArb_l261_1 = ({7'd0,1'b1} <<< fsm_rLkReq_0_wLen);
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_rLkReq_0_lkType)
      LkT_rd : fsm_rLkReq_0_lkType_string = "rd    ";
      LkT_wr : fsm_rLkReq_0_lkType_string = "wr    ";
      LkT_raw : fsm_rLkReq_0_lkType_string = "raw   ";
      LkT_insTab : fsm_rLkReq_0_lkType_string = "insTab";
      default : fsm_rLkReq_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_lkReqV_0_lkType)
      LkT_rd : fsm_lkReqV_0_lkType_string = "rd    ";
      LkT_wr : fsm_lkReqV_0_lkType_string = "wr    ";
      LkT_raw : fsm_lkReqV_0_lkType_string = "raw   ";
      LkT_insTab : fsm_lkReqV_0_lkType_string = "insTab";
      default : fsm_lkReqV_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_fsm_lkReqV_0_lkType)
      LkT_rd : _zz_fsm_lkReqV_0_lkType_string = "rd    ";
      LkT_wr : _zz_fsm_lkReqV_0_lkType_string = "wr    ";
      LkT_raw : _zz_fsm_lkReqV_0_lkType_string = "raw   ";
      LkT_insTab : _zz_fsm_lkReqV_0_lkType_string = "insTab";
      default : _zz_fsm_lkReqV_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_lkReq_payload_lkType)
      LkT_rd : _zz_io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_lkReq_payload_lkType_string = "insTab";
      default : _zz_io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_3_BOOT : fsm_stateReg_string = "BOOT     ";
      fsm_enumDef_3_LKREQ : fsm_stateReg_string = "LKREQ    ";
      fsm_enumDef_3_LKREQFIRE : fsm_stateReg_string = "LKREQFIRE";
      fsm_enumDef_3_WRDATA : fsm_stateReg_string = "WRDATA   ";
      default : fsm_stateReg_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_3_BOOT : fsm_stateNext_string = "BOOT     ";
      fsm_enumDef_3_LKREQ : fsm_stateNext_string = "LKREQ    ";
      fsm_enumDef_3_LKREQFIRE : fsm_stateNext_string = "LKREQFIRE";
      fsm_enumDef_3_WRDATA : fsm_stateNext_string = "WRDATA   ";
      default : fsm_stateNext_string = "?????????";
    endcase
  end
  `endif

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
      end
      fsm_enumDef_3_LKREQFIRE : begin
      end
      fsm_enumDef_3_WRDATA : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_cntFire_willIncrement = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
      end
      fsm_enumDef_3_LKREQFIRE : begin
        if(io_lkReq_fire) begin
          fsm_cntFire_willIncrement = 1'b1;
        end
      end
      fsm_enumDef_3_WRDATA : begin
      end
      default : begin
      end
    endcase
  end

  assign fsm_cntFire_willClear = 1'b0;
  assign fsm_cntFire_willOverflowIfInc = 1'b1;
  assign fsm_cntFire_willOverflow = (fsm_cntFire_willOverflowIfInc && fsm_cntFire_willIncrement);
  assign fsm_lkReqBitV_0 = _zz_fsm_lkReqBitV_0[46 : 0];
  assign fsm_lkReqV_0_nId = fsm_lkReqBitV_0[0 : 0];
  assign fsm_lkReqV_0_tId = fsm_lkReqBitV_0[22 : 1];
  assign fsm_lkReqV_0_tabId = fsm_lkReqBitV_0[25 : 23];
  assign fsm_lkReqV_0_snId = fsm_lkReqBitV_0[26 : 26];
  assign fsm_lkReqV_0_txnId = fsm_lkReqBitV_0[32 : 27];
  assign _zz_fsm_lkReqV_0_lkType = fsm_lkReqBitV_0[34 : 33];
  assign fsm_lkReqV_0_lkType = _zz_fsm_lkReqV_0_lkType;
  assign fsm_lkReqV_0_lkRelease = fsm_lkReqBitV_0[35];
  assign fsm_lkReqV_0_txnTimeOut = fsm_lkReqBitV_0[36];
  assign fsm_lkReqV_0_txnAbt = fsm_lkReqBitV_0[37];
  assign fsm_lkReqV_0_lkIdx = fsm_lkReqBitV_0[43 : 38];
  assign fsm_lkReqV_0_wLen = fsm_lkReqBitV_0[46 : 44];
  assign fsm_MskWr[0] = ((fsm_lkReqV_0_lkRelease && ((fsm_lkReqV_0_lkType == LkT_wr) || (fsm_lkReqV_0_lkType == LkT_raw))) && (! fsm_lkReqV_0_txnAbt));
  always @(*) begin
    io_lkReq_valid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
      end
      fsm_enumDef_3_LKREQFIRE : begin
        io_lkReq_valid = 1'b1;
      end
      fsm_enumDef_3_WRDATA : begin
      end
      default : begin
      end
    endcase
  end

  assign _zz_io_lkReq_payload_lkType = fsm_rLkReq_0_lkType;
  assign io_lkReq_payload_nId = fsm_rLkReq_0_nId;
  assign io_lkReq_payload_tId = fsm_rLkReq_0_tId;
  assign io_lkReq_payload_tabId = fsm_rLkReq_0_tabId;
  assign io_lkReq_payload_snId = fsm_rLkReq_0_snId;
  assign io_lkReq_payload_txnId = fsm_rLkReq_0_txnId;
  assign io_lkReq_payload_lkType = _zz_io_lkReq_payload_lkType;
  assign io_lkReq_payload_lkRelease = fsm_rLkReq_0_lkRelease;
  assign io_lkReq_payload_txnTimeOut = fsm_rLkReq_0_txnTimeOut;
  assign io_lkReq_payload_txnAbt = fsm_rLkReq_0_txnAbt;
  assign io_lkReq_payload_lkIdx = fsm_rLkReq_0_lkIdx;
  assign io_lkReq_payload_wLen = fsm_rLkReq_0_wLen;
  always @(*) begin
    io_reqQ_ready = (io_wrData_ready && _zz_io_reqQ_ready);
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
        io_reqQ_ready = 1'b1;
      end
      fsm_enumDef_3_LKREQFIRE : begin
      end
      fsm_enumDef_3_WRDATA : begin
        io_reqQ_ready = io_wrData_ready;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_wrData_valid = (io_reqQ_valid && _zz_io_reqQ_ready);
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
      end
      fsm_enumDef_3_LKREQFIRE : begin
      end
      fsm_enumDef_3_WRDATA : begin
        io_wrData_valid = io_reqQ_valid;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_wrData_payload = io_reqQ_payload;
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
      end
      fsm_enumDef_3_LKREQFIRE : begin
      end
      fsm_enumDef_3_WRDATA : begin
        io_wrData_payload = io_reqQ_payload;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
        if(io_reqQ_fire) begin
          fsm_stateNext = fsm_enumDef_3_LKREQFIRE;
        end
      end
      fsm_enumDef_3_LKREQFIRE : begin
        if(io_lkReq_fire) begin
          if(fsm_cntFire_willOverflow) begin
            case(switch_NetArb_l241)
              1'b1 : begin
                fsm_stateNext = fsm_enumDef_3_WRDATA;
              end
              default : begin
                fsm_stateNext = fsm_enumDef_3_LKREQ;
              end
            endcase
          end
        end
      end
      fsm_enumDef_3_WRDATA : begin
        if(io_reqQ_fire_1) begin
          if(when_NetArb_l261) begin
            if(when_NetArb_l265) begin
              fsm_stateNext = fsm_enumDef_3_LKREQ;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_3_LKREQ;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_3_BOOT;
    end
  end

  assign io_reqQ_fire = (io_reqQ_valid && io_reqQ_ready);
  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign switch_NetArb_l241 = (|fsm_rMskWr);
  assign fsm_rMskWr_ohFirst_input = fsm_rMskWr;
  assign fsm_rMskWr_ohFirst_masked = (fsm_rMskWr_ohFirst_input & (~ _zz_fsm_rMskWr_ohFirst_masked));
  assign fsm_rMskWr_ohFirst_value = fsm_rMskWr_ohFirst_masked;
  always @(*) begin
    _zz_when_NetArb_l265 = 1'b1;
    if(io_reqQ_fire_1) begin
      if(when_NetArb_l261) begin
        _zz_when_NetArb_l265[0] = 1'b0;
      end
    end
  end

  assign io_reqQ_fire_1 = (io_reqQ_valid && io_reqQ_ready);
  assign when_NetArb_l261 = (cntBeat == _zz_when_NetArb_l261);
  assign when_NetArb_l265 = (! (|(fsm_rMskWr & _zz_when_NetArb_l265)));
  assign _zz_io_reqQ_ready = (fsm_stateReg == fsm_enumDef_3_WRDATA);
  always @(posedge clk) begin
    if(!resetn) begin
      cntBeat <= 8'h0;
      fsm_rMskWr <= 1'b0;
      fsm_stateReg <= fsm_enumDef_3_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_3_LKREQ : begin
          if(io_reqQ_fire) begin
            fsm_rMskWr <= fsm_MskWr;
          end
        end
        fsm_enumDef_3_LKREQFIRE : begin
        end
        fsm_enumDef_3_WRDATA : begin
          if(io_reqQ_fire_1) begin
            cntBeat <= (cntBeat + 8'h01);
            if(when_NetArb_l261) begin
              fsm_rMskWr[0] <= 1'b0;
              cntBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_enumDef_3_LKREQ : begin
        if(io_reqQ_fire) begin
          fsm_rLkReq_0_nId <= fsm_lkReqV_0_nId;
          fsm_rLkReq_0_tId <= fsm_lkReqV_0_tId;
          fsm_rLkReq_0_tabId <= fsm_lkReqV_0_tabId;
          fsm_rLkReq_0_snId <= fsm_lkReqV_0_snId;
          fsm_rLkReq_0_txnId <= fsm_lkReqV_0_txnId;
          fsm_rLkReq_0_lkType <= fsm_lkReqV_0_lkType;
          fsm_rLkReq_0_lkRelease <= fsm_lkReqV_0_lkRelease;
          fsm_rLkReq_0_txnTimeOut <= fsm_lkReqV_0_txnTimeOut;
          fsm_rLkReq_0_txnAbt <= fsm_lkReqV_0_txnAbt;
          fsm_rLkReq_0_lkIdx <= fsm_lkReqV_0_lkIdx;
          fsm_rLkReq_0_wLen <= fsm_lkReqV_0_wLen;
        end
      end
      fsm_enumDef_3_LKREQFIRE : begin
      end
      fsm_enumDef_3_WRDATA : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module RecvDispatcher (
  input               io_recvQ_valid,
  output reg          io_recvQ_ready,
  input      [511:0]  io_recvQ_payload,
  output reg          io_lkRespV_0_valid,
  input               io_lkRespV_0_ready,
  output reg [0:0]    io_lkRespV_0_payload_nId,
  output reg [21:0]   io_lkRespV_0_payload_tId,
  output reg [2:0]    io_lkRespV_0_payload_tabId,
  output reg [0:0]    io_lkRespV_0_payload_snId,
  output reg [5:0]    io_lkRespV_0_payload_txnId,
  output reg [1:0]    io_lkRespV_0_payload_lkType,
  output reg          io_lkRespV_0_payload_lkRelease,
  output reg          io_lkRespV_0_payload_txnAbt,
  output reg [5:0]    io_lkRespV_0_payload_lkIdx,
  output reg [2:0]    io_lkRespV_0_payload_wLen,
  output reg [1:0]    io_lkRespV_0_payload_respType,
  output reg          io_lkRespV_0_payload_lkWaited,
  output reg          io_rdDataV_0_valid,
  input               io_rdDataV_0_ready,
  output reg [511:0]  io_rdDataV_0_payload,
  output              io_statusVld,
  output     [3:0]    io_nResp,
  output     [3:0]    io_nWrCmtResp,
  output     [3:0]    io_nRdGetResp,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam fsm_enumDef_2_BOOT = 2'd0;
  localparam fsm_enumDef_2_LKRESP = 2'd1;
  localparam fsm_enumDef_2_LKDISPATCH = 2'd2;
  localparam fsm_enumDef_2_RDDATA = 2'd3;

  wire       [48:0]   _zz_fsm_lkRespBitV_0;
  wire       [0:0]    _zz_io_nResp;
  reg        [0:0]    _zz_io_nWrCmtResp;
  wire       [0:0]    _zz_io_nWrCmtResp_1;
  reg        [0:0]    _zz_io_nRdGetResp;
  wire       [0:0]    _zz_io_nRdGetResp_1;
  wire       [0:0]    _zz__zz_1;
  wire                _zz_when;
  wire       [0:0]    _zz_fsm_rMskRd_ohFirst_masked;
  wire       [0:0]    _zz__zz_2;
  wire       [7:0]    _zz_when_NetArb_l173;
  wire       [7:0]    _zz_when_NetArb_l173_1;
  reg        [7:0]    cntBeat;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 fsm_cntDisp_willIncrement;
  wire                fsm_cntDisp_willClear;
  wire                fsm_cntDisp_willOverflowIfInc;
  wire                fsm_cntDisp_willOverflow;
  reg        [0:0]    fsm_rLkResp_0_nId;
  reg        [21:0]   fsm_rLkResp_0_tId;
  reg        [2:0]    fsm_rLkResp_0_tabId;
  reg        [0:0]    fsm_rLkResp_0_snId;
  reg        [5:0]    fsm_rLkResp_0_txnId;
  reg        [1:0]    fsm_rLkResp_0_lkType;
  reg                 fsm_rLkResp_0_lkRelease;
  reg                 fsm_rLkResp_0_txnAbt;
  reg        [5:0]    fsm_rLkResp_0_lkIdx;
  reg        [2:0]    fsm_rLkResp_0_wLen;
  reg        [1:0]    fsm_rLkResp_0_respType;
  reg                 fsm_rLkResp_0_lkWaited;
  wire       [48:0]   fsm_lkRespBitV_0;
  wire       [0:0]    fsm_lkRespV_0_nId;
  wire       [21:0]   fsm_lkRespV_0_tId;
  wire       [2:0]    fsm_lkRespV_0_tabId;
  wire       [0:0]    fsm_lkRespV_0_snId;
  wire       [5:0]    fsm_lkRespV_0_txnId;
  wire       [1:0]    fsm_lkRespV_0_lkType;
  wire                fsm_lkRespV_0_lkRelease;
  wire                fsm_lkRespV_0_txnAbt;
  wire       [5:0]    fsm_lkRespV_0_lkIdx;
  wire       [2:0]    fsm_lkRespV_0_wLen;
  wire       [1:0]    fsm_lkRespV_0_respType;
  wire                fsm_lkRespV_0_lkWaited;
  wire       [1:0]    _zz_fsm_lkRespV_0_lkType;
  wire       [1:0]    _zz_fsm_lkRespV_0_respType;
  reg        [0:0]    fsm_rMskRd;
  wire       [0:0]    fsm_mskRd;
  wire       [0:0]    fsm_mskRdResp;
  wire       [0:0]    fsm_mskWrCmt;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                io_recvQ_fire;
  wire       [1:0]    _zz_io_lkRespV_0_payload_lkType;
  wire       [1:0]    _zz_io_lkRespV_0_payload_respType;
  wire                _zz_1;
  wire                switch_NetArb_l153;
  wire       [0:0]    fsm_rMskRd_ohFirst_input;
  wire       [0:0]    fsm_rMskRd_ohFirst_masked;
  wire       [0:0]    fsm_rMskRd_ohFirst_value;
  reg        [0:0]    _zz_when_NetArb_l178;
  wire                _zz_2;
  wire                io_recvQ_fire_1;
  wire                when_NetArb_l173;
  wire                when_NetArb_l178;
  `ifndef SYNTHESIS
  reg [47:0] io_lkRespV_0_payload_lkType_string;
  reg [71:0] io_lkRespV_0_payload_respType_string;
  reg [47:0] fsm_rLkResp_0_lkType_string;
  reg [71:0] fsm_rLkResp_0_respType_string;
  reg [47:0] fsm_lkRespV_0_lkType_string;
  reg [71:0] fsm_lkRespV_0_respType_string;
  reg [47:0] _zz_fsm_lkRespV_0_lkType_string;
  reg [71:0] _zz_fsm_lkRespV_0_respType_string;
  reg [79:0] fsm_stateReg_string;
  reg [79:0] fsm_stateNext_string;
  reg [47:0] _zz_io_lkRespV_0_payload_lkType_string;
  reg [71:0] _zz_io_lkRespV_0_payload_respType_string;
  `endif


  assign _zz_when = (io_lkRespV_0_valid && io_lkRespV_0_ready);
  assign _zz_fsm_lkRespBitV_0 = io_recvQ_payload[48 : 0];
  assign _zz_io_nResp = 1'b1;
  assign _zz__zz_1 = 1'b1;
  assign _zz_fsm_rMskRd_ohFirst_masked = (fsm_rMskRd_ohFirst_input - 1'b1);
  assign _zz__zz_2 = 1'b1;
  assign _zz_when_NetArb_l173 = (_zz_when_NetArb_l173_1 - 8'h01);
  assign _zz_when_NetArb_l173_1 = ({7'd0,1'b1} <<< fsm_rLkResp_0_wLen);
  assign _zz_io_nWrCmtResp_1 = fsm_mskWrCmt[0];
  assign _zz_io_nRdGetResp_1 = fsm_mskRdResp[0];
  always @(*) begin
    case(_zz_io_nWrCmtResp_1)
      1'b0 : _zz_io_nWrCmtResp = 1'b0;
      default : _zz_io_nWrCmtResp = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_io_nRdGetResp_1)
      1'b0 : _zz_io_nRdGetResp = 1'b0;
      default : _zz_io_nRdGetResp = 1'b1;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkRespV_0_payload_lkType)
      LkT_rd : io_lkRespV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_lkRespV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_lkRespV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkRespV_0_payload_lkType_string = "insTab";
      default : io_lkRespV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkRespV_0_payload_respType)
      LockRespType_grant : io_lkRespV_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkRespV_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkRespV_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkRespV_0_payload_respType_string = "release_1";
      default : io_lkRespV_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_rLkResp_0_lkType)
      LkT_rd : fsm_rLkResp_0_lkType_string = "rd    ";
      LkT_wr : fsm_rLkResp_0_lkType_string = "wr    ";
      LkT_raw : fsm_rLkResp_0_lkType_string = "raw   ";
      LkT_insTab : fsm_rLkResp_0_lkType_string = "insTab";
      default : fsm_rLkResp_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_rLkResp_0_respType)
      LockRespType_grant : fsm_rLkResp_0_respType_string = "grant    ";
      LockRespType_abort : fsm_rLkResp_0_respType_string = "abort    ";
      LockRespType_waiting : fsm_rLkResp_0_respType_string = "waiting  ";
      LockRespType_release_1 : fsm_rLkResp_0_respType_string = "release_1";
      default : fsm_rLkResp_0_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_lkRespV_0_lkType)
      LkT_rd : fsm_lkRespV_0_lkType_string = "rd    ";
      LkT_wr : fsm_lkRespV_0_lkType_string = "wr    ";
      LkT_raw : fsm_lkRespV_0_lkType_string = "raw   ";
      LkT_insTab : fsm_lkRespV_0_lkType_string = "insTab";
      default : fsm_lkRespV_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_lkRespV_0_respType)
      LockRespType_grant : fsm_lkRespV_0_respType_string = "grant    ";
      LockRespType_abort : fsm_lkRespV_0_respType_string = "abort    ";
      LockRespType_waiting : fsm_lkRespV_0_respType_string = "waiting  ";
      LockRespType_release_1 : fsm_lkRespV_0_respType_string = "release_1";
      default : fsm_lkRespV_0_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_fsm_lkRespV_0_lkType)
      LkT_rd : _zz_fsm_lkRespV_0_lkType_string = "rd    ";
      LkT_wr : _zz_fsm_lkRespV_0_lkType_string = "wr    ";
      LkT_raw : _zz_fsm_lkRespV_0_lkType_string = "raw   ";
      LkT_insTab : _zz_fsm_lkRespV_0_lkType_string = "insTab";
      default : _zz_fsm_lkRespV_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_fsm_lkRespV_0_respType)
      LockRespType_grant : _zz_fsm_lkRespV_0_respType_string = "grant    ";
      LockRespType_abort : _zz_fsm_lkRespV_0_respType_string = "abort    ";
      LockRespType_waiting : _zz_fsm_lkRespV_0_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_fsm_lkRespV_0_respType_string = "release_1";
      default : _zz_fsm_lkRespV_0_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_2_BOOT : fsm_stateReg_string = "BOOT      ";
      fsm_enumDef_2_LKRESP : fsm_stateReg_string = "LKRESP    ";
      fsm_enumDef_2_LKDISPATCH : fsm_stateReg_string = "LKDISPATCH";
      fsm_enumDef_2_RDDATA : fsm_stateReg_string = "RDDATA    ";
      default : fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_2_BOOT : fsm_stateNext_string = "BOOT      ";
      fsm_enumDef_2_LKRESP : fsm_stateNext_string = "LKRESP    ";
      fsm_enumDef_2_LKDISPATCH : fsm_stateNext_string = "LKDISPATCH";
      fsm_enumDef_2_RDDATA : fsm_stateNext_string = "RDDATA    ";
      default : fsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_lkRespV_0_payload_lkType)
      LkT_rd : _zz_io_lkRespV_0_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_lkRespV_0_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_lkRespV_0_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_lkRespV_0_payload_lkType_string = "insTab";
      default : _zz_io_lkRespV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_lkRespV_0_payload_respType)
      LockRespType_grant : _zz_io_lkRespV_0_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_io_lkRespV_0_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_io_lkRespV_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_io_lkRespV_0_payload_respType_string = "release_1";
      default : _zz_io_lkRespV_0_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    fsm_cntDisp_willIncrement = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_when) begin
          fsm_cntDisp_willIncrement = 1'b1;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  assign fsm_cntDisp_willClear = 1'b0;
  assign fsm_cntDisp_willOverflowIfInc = 1'b1;
  assign fsm_cntDisp_willOverflow = (fsm_cntDisp_willOverflowIfInc && fsm_cntDisp_willIncrement);
  assign fsm_lkRespBitV_0 = _zz_fsm_lkRespBitV_0[48 : 0];
  assign fsm_lkRespV_0_nId = fsm_lkRespBitV_0[0 : 0];
  assign fsm_lkRespV_0_tId = fsm_lkRespBitV_0[22 : 1];
  assign fsm_lkRespV_0_tabId = fsm_lkRespBitV_0[25 : 23];
  assign fsm_lkRespV_0_snId = fsm_lkRespBitV_0[26 : 26];
  assign fsm_lkRespV_0_txnId = fsm_lkRespBitV_0[32 : 27];
  assign _zz_fsm_lkRespV_0_lkType = fsm_lkRespBitV_0[34 : 33];
  assign fsm_lkRespV_0_lkType = _zz_fsm_lkRespV_0_lkType;
  assign fsm_lkRespV_0_lkRelease = fsm_lkRespBitV_0[35];
  assign fsm_lkRespV_0_txnAbt = fsm_lkRespBitV_0[36];
  assign fsm_lkRespV_0_lkIdx = fsm_lkRespBitV_0[42 : 37];
  assign fsm_lkRespV_0_wLen = fsm_lkRespBitV_0[45 : 43];
  assign _zz_fsm_lkRespV_0_respType = fsm_lkRespBitV_0[47 : 46];
  assign fsm_lkRespV_0_respType = _zz_fsm_lkRespV_0_respType;
  assign fsm_lkRespV_0_lkWaited = fsm_lkRespBitV_0[48];
  assign fsm_mskRd[0] = (((! fsm_lkRespV_0_lkRelease) && ((fsm_lkRespV_0_lkType == LkT_rd) || (fsm_lkRespV_0_lkType == LkT_raw))) && (fsm_lkRespV_0_respType == LockRespType_grant));
  assign fsm_mskRdResp[0] = ((! fsm_lkRespV_0_lkRelease) && ((fsm_lkRespV_0_lkType == LkT_rd) || (fsm_lkRespV_0_lkType == LkT_raw)));
  assign fsm_mskWrCmt[0] = ((fsm_lkRespV_0_lkRelease && ((fsm_lkRespV_0_lkType == LkT_wr) || (fsm_lkRespV_0_lkType == LkT_raw))) && (! fsm_lkRespV_0_txnAbt));
  always @(*) begin
    io_recvQ_ready = (fsm_stateReg == fsm_enumDef_2_LKRESP);
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
      end
      fsm_enumDef_2_RDDATA : begin
        io_recvQ_ready = io_rdDataV_0_ready;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_valid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_valid = 1'b1;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_nId = 1'bx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_nId = fsm_rLkResp_0_nId;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_tId = 22'bxxxxxxxxxxxxxxxxxxxxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_tId = fsm_rLkResp_0_tId;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_tabId = 3'bxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_tabId = fsm_rLkResp_0_tabId;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_snId = 1'bx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_snId = fsm_rLkResp_0_snId;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_txnId = 6'bxxxxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_txnId = fsm_rLkResp_0_txnId;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_lkType = (2'bxx);
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_lkType = _zz_io_lkRespV_0_payload_lkType;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_lkRelease = 1'bx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_lkRelease = fsm_rLkResp_0_lkRelease;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_txnAbt = 1'bx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_txnAbt = fsm_rLkResp_0_txnAbt;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_lkIdx = 6'bxxxxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_lkIdx = fsm_rLkResp_0_lkIdx;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_wLen = 3'bxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_wLen = fsm_rLkResp_0_wLen;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_respType = (2'bxx);
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_respType = _zz_io_lkRespV_0_payload_respType;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkRespV_0_payload_lkWaited = 1'bx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_1) begin
          io_lkRespV_0_payload_lkWaited = fsm_rLkResp_0_lkWaited;
        end
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_rdDataV_0_valid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
      end
      fsm_enumDef_2_RDDATA : begin
        if(_zz_2) begin
          io_rdDataV_0_valid = io_recvQ_valid;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_rdDataV_0_payload = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
      end
      fsm_enumDef_2_LKDISPATCH : begin
      end
      fsm_enumDef_2_RDDATA : begin
        if(_zz_2) begin
          io_rdDataV_0_payload = io_recvQ_payload;
        end
      end
      default : begin
      end
    endcase
  end

  assign io_statusVld = (fsm_stateReg == fsm_enumDef_2_LKRESP);
  assign io_nResp = {3'd0, _zz_io_nResp};
  assign io_nWrCmtResp = {3'd0, _zz_io_nWrCmtResp};
  assign io_nRdGetResp = {3'd0, _zz_io_nRdGetResp};
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
        if(io_recvQ_fire) begin
          fsm_stateNext = fsm_enumDef_2_LKDISPATCH;
        end
      end
      fsm_enumDef_2_LKDISPATCH : begin
        if(_zz_when) begin
          if(fsm_cntDisp_willOverflow) begin
            case(switch_NetArb_l153)
              1'b1 : begin
                fsm_stateNext = fsm_enumDef_2_RDDATA;
              end
              default : begin
                fsm_stateNext = fsm_enumDef_2_LKRESP;
              end
            endcase
          end
        end
      end
      fsm_enumDef_2_RDDATA : begin
        if(io_recvQ_fire_1) begin
          if(when_NetArb_l173) begin
            if(when_NetArb_l178) begin
              fsm_stateNext = fsm_enumDef_2_LKRESP;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_2_LKRESP;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_2_BOOT;
    end
  end

  assign io_recvQ_fire = (io_recvQ_valid && io_recvQ_ready);
  assign _zz_io_lkRespV_0_payload_lkType = fsm_rLkResp_0_lkType;
  assign _zz_io_lkRespV_0_payload_respType = fsm_rLkResp_0_respType;
  assign _zz_1 = _zz__zz_1[0];
  assign switch_NetArb_l153 = (|fsm_rMskRd);
  assign fsm_rMskRd_ohFirst_input = fsm_rMskRd;
  assign fsm_rMskRd_ohFirst_masked = (fsm_rMskRd_ohFirst_input & (~ _zz_fsm_rMskRd_ohFirst_masked));
  assign fsm_rMskRd_ohFirst_value = fsm_rMskRd_ohFirst_masked;
  always @(*) begin
    _zz_when_NetArb_l178 = 1'b1;
    if(io_recvQ_fire_1) begin
      if(when_NetArb_l173) begin
        _zz_when_NetArb_l178[0] = 1'b0;
      end
    end
  end

  assign _zz_2 = _zz__zz_2[0];
  assign io_recvQ_fire_1 = (io_recvQ_valid && io_recvQ_ready);
  assign when_NetArb_l173 = (cntBeat == _zz_when_NetArb_l173);
  assign when_NetArb_l178 = (! (|(fsm_rMskRd & _zz_when_NetArb_l178)));
  always @(posedge clk) begin
    if(!resetn) begin
      cntBeat <= 8'h0;
      fsm_rMskRd <= 1'b0;
      fsm_stateReg <= fsm_enumDef_2_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_2_LKRESP : begin
          if(io_recvQ_fire) begin
            fsm_rMskRd <= fsm_mskRd;
          end
        end
        fsm_enumDef_2_LKDISPATCH : begin
        end
        fsm_enumDef_2_RDDATA : begin
          if(io_recvQ_fire_1) begin
            cntBeat <= (cntBeat + 8'h01);
            if(when_NetArb_l173) begin
              fsm_rMskRd[0] <= 1'b0;
              cntBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_enumDef_2_LKRESP : begin
        if(io_recvQ_fire) begin
          fsm_rLkResp_0_nId <= fsm_lkRespV_0_nId;
          fsm_rLkResp_0_tId <= fsm_lkRespV_0_tId;
          fsm_rLkResp_0_tabId <= fsm_lkRespV_0_tabId;
          fsm_rLkResp_0_snId <= fsm_lkRespV_0_snId;
          fsm_rLkResp_0_txnId <= fsm_lkRespV_0_txnId;
          fsm_rLkResp_0_lkType <= fsm_lkRespV_0_lkType;
          fsm_rLkResp_0_lkRelease <= fsm_lkRespV_0_lkRelease;
          fsm_rLkResp_0_txnAbt <= fsm_lkRespV_0_txnAbt;
          fsm_rLkResp_0_lkIdx <= fsm_lkRespV_0_lkIdx;
          fsm_rLkResp_0_wLen <= fsm_lkRespV_0_wLen;
          fsm_rLkResp_0_respType <= fsm_lkRespV_0_respType;
          fsm_rLkResp_0_lkWaited <= fsm_lkRespV_0_lkWaited;
        end
      end
      fsm_enumDef_2_LKDISPATCH : begin
      end
      fsm_enumDef_2_RDDATA : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module SendArbiter (
  input               io_lkReqV_0_valid,
  output              io_lkReqV_0_ready,
  input      [0:0]    io_lkReqV_0_payload_nId,
  input      [21:0]   io_lkReqV_0_payload_tId,
  input      [2:0]    io_lkReqV_0_payload_tabId,
  input      [0:0]    io_lkReqV_0_payload_snId,
  input      [5:0]    io_lkReqV_0_payload_txnId,
  input      [1:0]    io_lkReqV_0_payload_lkType,
  input               io_lkReqV_0_payload_lkRelease,
  input               io_lkReqV_0_payload_txnTimeOut,
  input               io_lkReqV_0_payload_txnAbt,
  input      [5:0]    io_lkReqV_0_payload_lkIdx,
  input      [2:0]    io_lkReqV_0_payload_wLen,
  input               io_wrDataV_0_valid,
  output reg          io_wrDataV_0_ready,
  input      [511:0]  io_wrDataV_0_payload,
  output reg          io_sendQ_valid,
  input               io_sendQ_ready,
  output reg [511:0]  io_sendQ_payload,
  output              io_statusVld,
  output     [3:0]    io_nReq,
  output     [3:0]    io_nWrCmtReq,
  output     [3:0]    io_nRdGetReq,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam fsm_enumDef_1_BOOT = 2'd0;
  localparam fsm_enumDef_1_LKREQ = 2'd1;
  localparam fsm_enumDef_1_WRDATA = 2'd2;

  wire       [46:0]   _zz_lkReqJoin_payload;
  wire       [0:0]    _zz_io_nReq;
  reg        [0:0]    _zz_io_nWrCmtReq;
  wire       [0:0]    _zz_io_nWrCmtReq_1;
  reg        [0:0]    _zz_io_nRdGetReq;
  wire       [0:0]    _zz_io_nRdGetReq_1;
  wire       [0:0]    _zz_fsm_rMskWr_ohFirst_masked;
  wire       [0:0]    _zz_when;
  wire       [7:0]    _zz_when_NetArb_l75;
  wire       [7:0]    _zz_when_NetArb_l75_1;
  wire                lkReqJoin_valid;
  wire                lkReqJoin_ready;
  wire       [511:0]  lkReqJoin_payload;
  wire                tmpJoin_valid;
  wire                tmpJoin_ready;
  wire       [0:0]    tmpJoin_payload_0_nId;
  wire       [21:0]   tmpJoin_payload_0_tId;
  wire       [2:0]    tmpJoin_payload_0_tabId;
  wire       [0:0]    tmpJoin_payload_0_snId;
  wire       [5:0]    tmpJoin_payload_0_txnId;
  wire       [1:0]    tmpJoin_payload_0_lkType;
  wire                tmpJoin_payload_0_lkRelease;
  wire                tmpJoin_payload_0_txnTimeOut;
  wire                tmpJoin_payload_0_txnAbt;
  wire       [5:0]    tmpJoin_payload_0_lkIdx;
  wire       [2:0]    tmpJoin_payload_0_wLen;
  wire                tmpJoin_fire;
  reg        [2:0]    rWrLen_0;
  reg        [7:0]    cntBeat;
  wire       [0:0]    mskWr;
  wire       [0:0]    mskRdGet;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [0:0]    fsm_rMskWr;
  wire                _zz_io_sendQ_valid;
  reg        [1:0]    fsm_stateReg;
  reg        [1:0]    fsm_stateNext;
  wire                io_sendQ_fire;
  wire                when_NetArb_l59;
  wire       [0:0]    fsm_rMskWr_ohFirst_input;
  wire       [0:0]    fsm_rMskWr_ohFirst_masked;
  wire       [0:0]    fsm_rMskWr_ohFirst_value;
  reg        [0:0]    _zz_when_NetArb_l80;
  wire                io_sendQ_fire_1;
  wire                when_NetArb_l75;
  wire                when_NetArb_l80;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReqV_0_payload_lkType_string;
  reg [47:0] tmpJoin_payload_0_lkType_string;
  reg [47:0] fsm_stateReg_string;
  reg [47:0] fsm_stateNext_string;
  `endif


  assign _zz_lkReqJoin_payload = {tmpJoin_payload_0_wLen,{tmpJoin_payload_0_lkIdx,{tmpJoin_payload_0_txnAbt,{tmpJoin_payload_0_txnTimeOut,{tmpJoin_payload_0_lkRelease,{tmpJoin_payload_0_lkType,{tmpJoin_payload_0_txnId,{tmpJoin_payload_0_snId,{tmpJoin_payload_0_tabId,{tmpJoin_payload_0_tId,tmpJoin_payload_0_nId}}}}}}}}}};
  assign _zz_io_nReq = 1'b1;
  assign _zz_fsm_rMskWr_ohFirst_masked = (fsm_rMskWr_ohFirst_input - 1'b1);
  assign _zz_when = 1'b1;
  assign _zz_when_NetArb_l75 = (_zz_when_NetArb_l75_1 - 8'h01);
  assign _zz_when_NetArb_l75_1 = ({7'd0,1'b1} <<< rWrLen_0);
  assign _zz_io_nWrCmtReq_1 = mskWr[0];
  assign _zz_io_nRdGetReq_1 = mskRdGet[0];
  always @(*) begin
    case(_zz_io_nWrCmtReq_1)
      1'b0 : _zz_io_nWrCmtReq = 1'b0;
      default : _zz_io_nWrCmtReq = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_io_nRdGetReq_1)
      1'b0 : _zz_io_nRdGetReq = 1'b0;
      default : _zz_io_nRdGetReq = 1'b1;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReqV_0_payload_lkType)
      LkT_rd : io_lkReqV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReqV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReqV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReqV_0_payload_lkType_string = "insTab";
      default : io_lkReqV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(tmpJoin_payload_0_lkType)
      LkT_rd : tmpJoin_payload_0_lkType_string = "rd    ";
      LkT_wr : tmpJoin_payload_0_lkType_string = "wr    ";
      LkT_raw : tmpJoin_payload_0_lkType_string = "raw   ";
      LkT_insTab : tmpJoin_payload_0_lkType_string = "insTab";
      default : tmpJoin_payload_0_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_1_BOOT : fsm_stateReg_string = "BOOT  ";
      fsm_enumDef_1_LKREQ : fsm_stateReg_string = "LKREQ ";
      fsm_enumDef_1_WRDATA : fsm_stateReg_string = "WRDATA";
      default : fsm_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_1_BOOT : fsm_stateNext_string = "BOOT  ";
      fsm_enumDef_1_LKREQ : fsm_stateNext_string = "LKREQ ";
      fsm_enumDef_1_WRDATA : fsm_stateNext_string = "WRDATA";
      default : fsm_stateNext_string = "??????";
    endcase
  end
  `endif

  assign tmpJoin_payload_0_nId = io_lkReqV_0_payload_nId;
  assign tmpJoin_payload_0_tId = io_lkReqV_0_payload_tId;
  assign tmpJoin_payload_0_tabId = io_lkReqV_0_payload_tabId;
  assign tmpJoin_payload_0_snId = io_lkReqV_0_payload_snId;
  assign tmpJoin_payload_0_txnId = io_lkReqV_0_payload_txnId;
  assign tmpJoin_payload_0_lkType = io_lkReqV_0_payload_lkType;
  assign tmpJoin_payload_0_lkRelease = io_lkReqV_0_payload_lkRelease;
  assign tmpJoin_payload_0_txnTimeOut = io_lkReqV_0_payload_txnTimeOut;
  assign tmpJoin_payload_0_txnAbt = io_lkReqV_0_payload_txnAbt;
  assign tmpJoin_payload_0_lkIdx = io_lkReqV_0_payload_lkIdx;
  assign tmpJoin_payload_0_wLen = io_lkReqV_0_payload_wLen;
  assign tmpJoin_valid = io_lkReqV_0_valid;
  assign tmpJoin_fire = (tmpJoin_valid && tmpJoin_ready);
  assign io_lkReqV_0_ready = tmpJoin_fire;
  assign lkReqJoin_valid = tmpJoin_valid;
  assign tmpJoin_ready = lkReqJoin_ready;
  assign lkReqJoin_payload = {465'd0, _zz_lkReqJoin_payload};
  assign mskWr[0] = ((io_lkReqV_0_payload_lkRelease && ((io_lkReqV_0_payload_lkType == LkT_wr) || (io_lkReqV_0_payload_lkType == LkT_raw))) && (! io_lkReqV_0_payload_txnAbt));
  assign mskRdGet[0] = ((! io_lkReqV_0_payload_lkRelease) && ((io_lkReqV_0_payload_lkType == LkT_rd) || (io_lkReqV_0_payload_lkType == LkT_raw)));
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
      end
      fsm_enumDef_1_WRDATA : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    io_wrDataV_0_ready = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
      end
      fsm_enumDef_1_WRDATA : begin
        if(_zz_when[0]) begin
          io_wrDataV_0_ready = io_sendQ_ready;
        end
      end
      default : begin
      end
    endcase
  end

  assign lkReqJoin_ready = (io_sendQ_ready && _zz_io_sendQ_valid);
  always @(*) begin
    io_sendQ_valid = (lkReqJoin_valid && _zz_io_sendQ_valid);
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
      end
      fsm_enumDef_1_WRDATA : begin
        io_sendQ_valid = io_wrDataV_0_valid;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_sendQ_payload = lkReqJoin_payload;
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
      end
      fsm_enumDef_1_WRDATA : begin
        io_sendQ_payload = io_wrDataV_0_payload;
      end
      default : begin
      end
    endcase
  end

  assign io_statusVld = (fsm_stateReg == fsm_enumDef_1_LKREQ);
  assign io_nReq = {3'd0, _zz_io_nReq};
  assign io_nWrCmtReq = {3'd0, _zz_io_nWrCmtReq};
  assign io_nRdGetReq = {3'd0, _zz_io_nRdGetReq};
  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
        if(io_sendQ_fire) begin
          if(when_NetArb_l59) begin
            fsm_stateNext = fsm_enumDef_1_WRDATA;
          end
        end
      end
      fsm_enumDef_1_WRDATA : begin
        if(io_sendQ_fire_1) begin
          if(when_NetArb_l75) begin
            if(when_NetArb_l80) begin
              fsm_stateNext = fsm_enumDef_1_LKREQ;
            end
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_1_LKREQ;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_1_BOOT;
    end
  end

  assign io_sendQ_fire = (io_sendQ_valid && io_sendQ_ready);
  assign when_NetArb_l59 = (|mskWr);
  assign fsm_rMskWr_ohFirst_input = fsm_rMskWr;
  assign fsm_rMskWr_ohFirst_masked = (fsm_rMskWr_ohFirst_input & (~ _zz_fsm_rMskWr_ohFirst_masked));
  assign fsm_rMskWr_ohFirst_value = fsm_rMskWr_ohFirst_masked;
  always @(*) begin
    _zz_when_NetArb_l80 = 1'b1;
    if(io_sendQ_fire_1) begin
      if(when_NetArb_l75) begin
        _zz_when_NetArb_l80[0] = 1'b0;
      end
    end
  end

  assign io_sendQ_fire_1 = (io_sendQ_valid && io_sendQ_ready);
  assign when_NetArb_l75 = (cntBeat == _zz_when_NetArb_l75);
  assign when_NetArb_l80 = (! (|(fsm_rMskWr & _zz_when_NetArb_l80)));
  assign _zz_io_sendQ_valid = (fsm_stateReg == fsm_enumDef_1_LKREQ);
  always @(posedge clk) begin
    if(!resetn) begin
      cntBeat <= 8'h0;
      fsm_rMskWr <= 1'b0;
      fsm_stateReg <= fsm_enumDef_1_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_1_LKREQ : begin
          if(io_sendQ_fire) begin
            fsm_rMskWr <= mskWr;
          end
        end
        fsm_enumDef_1_WRDATA : begin
          if(io_sendQ_fire_1) begin
            cntBeat <= (cntBeat + 8'h01);
            if(when_NetArb_l75) begin
              fsm_rMskWr[0] <= 1'b0;
              cntBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_enumDef_1_LKREQ : begin
        if(io_sendQ_fire) begin
          rWrLen_0 <= io_lkReqV_0_payload_wLen;
        end
      end
      fsm_enumDef_1_WRDATA : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module TxnAgent (
  input               io_lkReq_valid,
  output              io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [21:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  input               io_wrData_valid,
  output              io_wrData_ready,
  input      [511:0]  io_wrData_payload,
  output reg          io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [21:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  output              io_rdData_valid,
  input               io_rdData_ready,
  output     [511:0]  io_rdData_payload,
  output              io_axi_aw_valid,
  input               io_axi_aw_ready,
  output     [63:0]   io_axi_aw_payload_addr,
  output     [5:0]    io_axi_aw_payload_id,
  output     [7:0]    io_axi_aw_payload_len,
  output     [2:0]    io_axi_aw_payload_size,
  output     [1:0]    io_axi_aw_payload_burst,
  output              io_axi_w_valid,
  input               io_axi_w_ready,
  output     [511:0]  io_axi_w_payload_data,
  output     [63:0]   io_axi_w_payload_strb,
  output              io_axi_w_payload_last,
  input               io_axi_b_valid,
  output              io_axi_b_ready,
  input      [5:0]    io_axi_b_payload_id,
  input      [1:0]    io_axi_b_payload_resp,
  output reg          io_axi_ar_valid,
  input               io_axi_ar_ready,
  output     [63:0]   io_axi_ar_payload_addr,
  output     [5:0]    io_axi_ar_payload_id,
  output     [7:0]    io_axi_ar_payload_len,
  output     [2:0]    io_axi_ar_payload_size,
  output     [1:0]    io_axi_ar_payload_burst,
  input               io_axi_r_valid,
  output              io_axi_r_ready,
  input      [511:0]  io_axi_r_payload_data,
  input      [5:0]    io_axi_r_payload_id,
  input      [1:0]    io_axi_r_payload_resp,
  input               io_axi_r_payload_last,
  output              io_ltReq_valid,
  input               io_ltReq_ready,
  output     [0:0]    io_ltReq_payload_nId,
  output     [21:0]   io_ltReq_payload_tId,
  output     [2:0]    io_ltReq_payload_tabId,
  output     [0:0]    io_ltReq_payload_snId,
  output     [5:0]    io_ltReq_payload_txnId,
  output     [1:0]    io_ltReq_payload_lkType,
  output              io_ltReq_payload_lkRelease,
  output              io_ltReq_payload_txnTimeOut,
  output              io_ltReq_payload_txnAbt,
  output     [5:0]    io_ltReq_payload_lkIdx,
  output     [2:0]    io_ltReq_payload_wLen,
  input               io_ltResp_valid,
  output reg          io_ltResp_ready,
  input      [0:0]    io_ltResp_payload_nId,
  input      [21:0]   io_ltResp_payload_tId,
  input      [2:0]    io_ltResp_payload_tabId,
  input      [0:0]    io_ltResp_payload_snId,
  input      [5:0]    io_ltResp_payload_txnId,
  input      [1:0]    io_ltResp_payload_lkType,
  input               io_ltResp_payload_lkRelease,
  input               io_ltResp_payload_txnAbt,
  input      [5:0]    io_ltResp_payload_lkIdx,
  input      [2:0]    io_ltResp_payload_wLen,
  input      [1:0]    io_ltResp_payload_respType,
  input               io_ltResp_payload_lkWaited,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                lkReqRlseWrFifo_io_pop_ready;
  wire       [0:0]    streamDemux_7_io_select;
  wire                streamArbiter_8_io_inputs_1_valid;
  wire       [2:0]    nBeatQ_io_push_payload;
  wire                nBeatQ_io_pop_ready;
  wire                io_lkReq_fifo_io_push_ready;
  wire                io_lkReq_fifo_io_pop_valid;
  wire       [0:0]    io_lkReq_fifo_io_pop_payload_nId;
  wire       [21:0]   io_lkReq_fifo_io_pop_payload_tId;
  wire       [2:0]    io_lkReq_fifo_io_pop_payload_tabId;
  wire       [0:0]    io_lkReq_fifo_io_pop_payload_snId;
  wire       [5:0]    io_lkReq_fifo_io_pop_payload_txnId;
  wire       [1:0]    io_lkReq_fifo_io_pop_payload_lkType;
  wire                io_lkReq_fifo_io_pop_payload_lkRelease;
  wire                io_lkReq_fifo_io_pop_payload_txnTimeOut;
  wire                io_lkReq_fifo_io_pop_payload_txnAbt;
  wire       [5:0]    io_lkReq_fifo_io_pop_payload_lkIdx;
  wire       [2:0]    io_lkReq_fifo_io_pop_payload_wLen;
  wire       [3:0]    io_lkReq_fifo_io_occupancy;
  wire       [3:0]    io_lkReq_fifo_io_availability;
  wire                lkReqRlseWrFifo_io_push_ready;
  wire                lkReqRlseWrFifo_io_pop_valid;
  wire       [0:0]    lkReqRlseWrFifo_io_pop_payload_nId;
  wire       [21:0]   lkReqRlseWrFifo_io_pop_payload_tId;
  wire       [2:0]    lkReqRlseWrFifo_io_pop_payload_tabId;
  wire       [0:0]    lkReqRlseWrFifo_io_pop_payload_snId;
  wire       [5:0]    lkReqRlseWrFifo_io_pop_payload_txnId;
  wire       [1:0]    lkReqRlseWrFifo_io_pop_payload_lkType;
  wire                lkReqRlseWrFifo_io_pop_payload_lkRelease;
  wire                lkReqRlseWrFifo_io_pop_payload_txnTimeOut;
  wire                lkReqRlseWrFifo_io_pop_payload_txnAbt;
  wire       [5:0]    lkReqRlseWrFifo_io_pop_payload_lkIdx;
  wire       [2:0]    lkReqRlseWrFifo_io_pop_payload_wLen;
  wire       [3:0]    lkReqRlseWrFifo_io_occupancy;
  wire       [3:0]    lkReqRlseWrFifo_io_availability;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [0:0]    streamDemux_7_io_outputs_0_payload_nId;
  wire       [21:0]   streamDemux_7_io_outputs_0_payload_tId;
  wire       [2:0]    streamDemux_7_io_outputs_0_payload_tabId;
  wire       [0:0]    streamDemux_7_io_outputs_0_payload_snId;
  wire       [5:0]    streamDemux_7_io_outputs_0_payload_txnId;
  wire       [1:0]    streamDemux_7_io_outputs_0_payload_lkType;
  wire                streamDemux_7_io_outputs_0_payload_lkRelease;
  wire                streamDemux_7_io_outputs_0_payload_txnTimeOut;
  wire                streamDemux_7_io_outputs_0_payload_txnAbt;
  wire       [5:0]    streamDemux_7_io_outputs_0_payload_lkIdx;
  wire       [2:0]    streamDemux_7_io_outputs_0_payload_wLen;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [0:0]    streamDemux_7_io_outputs_1_payload_nId;
  wire       [21:0]   streamDemux_7_io_outputs_1_payload_tId;
  wire       [2:0]    streamDemux_7_io_outputs_1_payload_tabId;
  wire       [0:0]    streamDemux_7_io_outputs_1_payload_snId;
  wire       [5:0]    streamDemux_7_io_outputs_1_payload_txnId;
  wire       [1:0]    streamDemux_7_io_outputs_1_payload_lkType;
  wire                streamDemux_7_io_outputs_1_payload_lkRelease;
  wire                streamDemux_7_io_outputs_1_payload_txnTimeOut;
  wire                streamDemux_7_io_outputs_1_payload_txnAbt;
  wire       [5:0]    streamDemux_7_io_outputs_1_payload_lkIdx;
  wire       [2:0]    streamDemux_7_io_outputs_1_payload_wLen;
  wire                streamArbiter_8_io_inputs_0_ready;
  wire                streamArbiter_8_io_inputs_1_ready;
  wire                streamArbiter_8_io_output_valid;
  wire       [0:0]    streamArbiter_8_io_output_payload_nId;
  wire       [21:0]   streamArbiter_8_io_output_payload_tId;
  wire       [2:0]    streamArbiter_8_io_output_payload_tabId;
  wire       [0:0]    streamArbiter_8_io_output_payload_snId;
  wire       [5:0]    streamArbiter_8_io_output_payload_txnId;
  wire       [1:0]    streamArbiter_8_io_output_payload_lkType;
  wire                streamArbiter_8_io_output_payload_lkRelease;
  wire                streamArbiter_8_io_output_payload_txnTimeOut;
  wire                streamArbiter_8_io_output_payload_txnAbt;
  wire       [5:0]    streamArbiter_8_io_output_payload_lkIdx;
  wire       [2:0]    streamArbiter_8_io_output_payload_wLen;
  wire       [0:0]    streamArbiter_8_io_chosen;
  wire       [1:0]    streamArbiter_8_io_chosenOH;
  wire                nBeatQ_io_push_ready;
  wire                nBeatQ_io_pop_valid;
  wire       [2:0]    nBeatQ_io_pop_payload;
  wire       [3:0]    nBeatQ_io_occupancy;
  wire                io_wrData_fifo_io_push_ready;
  wire                io_wrData_fifo_io_pop_valid;
  wire       [511:0]  io_wrData_fifo_io_pop_payload;
  wire       [3:0]    io_wrData_fifo_io_occupancy;
  wire       [3:0]    io_wrData_fifo_io_availability;
  wire       [27:0]   _zz_io_axi_aw_payload_addr;
  wire       [27:0]   _zz_io_axi_aw_payload_addr_1;
  wire       [7:0]    _zz_io_axi_aw_payload_len;
  wire       [7:0]    _zz_io_push_payload;
  wire       [7:0]    _zz_io_push_payload_1;
  wire       [2:0]    _zz_cntBeat_valueNext;
  wire       [0:0]    _zz_cntBeat_valueNext_1;
  wire       [27:0]   _zz_io_axi_ar_payload_addr;
  wire       [27:0]   _zz_io_axi_ar_payload_addr_1;
  wire       [7:0]    _zz_io_axi_ar_payload_len;
  wire                isWrReqRlse;
  wire                lkReqQFork_valid;
  reg                 lkReqQFork_ready;
  wire       [0:0]    lkReqQFork_payload_nId;
  wire       [21:0]   lkReqQFork_payload_tId;
  wire       [2:0]    lkReqQFork_payload_tabId;
  wire       [0:0]    lkReqQFork_payload_snId;
  wire       [5:0]    lkReqQFork_payload_txnId;
  wire       [1:0]    lkReqQFork_payload_lkType;
  wire                lkReqQFork_payload_lkRelease;
  wire                lkReqQFork_payload_txnTimeOut;
  wire                lkReqQFork_payload_txnAbt;
  wire       [5:0]    lkReqQFork_payload_lkIdx;
  wire       [2:0]    lkReqQFork_payload_wLen;
  wire                lkReqBpss_valid;
  wire                lkReqBpss_ready;
  wire       [0:0]    lkReqBpss_payload_nId;
  wire       [21:0]   lkReqBpss_payload_tId;
  wire       [2:0]    lkReqBpss_payload_tabId;
  wire       [0:0]    lkReqBpss_payload_snId;
  wire       [5:0]    lkReqBpss_payload_txnId;
  wire       [1:0]    lkReqBpss_payload_lkType;
  wire                lkReqBpss_payload_lkRelease;
  wire                lkReqBpss_payload_txnTimeOut;
  wire                lkReqBpss_payload_txnAbt;
  wire       [5:0]    lkReqBpss_payload_lkIdx;
  wire       [2:0]    lkReqBpss_payload_wLen;
  wire                io_axi_b_fire;
  reg        [3:0]    _zz_io_pop_ready;
  wire                lkReqRlseWrFifo_io_pop_fire;
  wire       [1:0]    switch_Helpers_l20;
  wire                _zz_io_pop_ready_1;
  wire       [1:0]    _zz_io_inputs_1_payload_lkType;
  wire                reqFork1_valid;
  wire                reqFork1_ready;
  wire       [0:0]    reqFork1_payload_nId;
  wire       [21:0]   reqFork1_payload_tId;
  wire       [2:0]    reqFork1_payload_tabId;
  wire       [0:0]    reqFork1_payload_snId;
  wire       [5:0]    reqFork1_payload_txnId;
  wire       [1:0]    reqFork1_payload_lkType;
  wire                reqFork1_payload_lkRelease;
  wire                reqFork1_payload_txnTimeOut;
  wire                reqFork1_payload_txnAbt;
  wire       [5:0]    reqFork1_payload_lkIdx;
  wire       [2:0]    reqFork1_payload_wLen;
  wire                reqFork2_valid;
  wire                reqFork2_ready;
  wire       [0:0]    reqFork2_payload_nId;
  wire       [21:0]   reqFork2_payload_tId;
  wire       [2:0]    reqFork2_payload_tabId;
  wire       [0:0]    reqFork2_payload_snId;
  wire       [5:0]    reqFork2_payload_txnId;
  wire       [1:0]    reqFork2_payload_lkType;
  wire                reqFork2_payload_lkRelease;
  wire                reqFork2_payload_txnTimeOut;
  wire                reqFork2_payload_txnAbt;
  wire       [5:0]    reqFork2_payload_lkIdx;
  wire       [2:0]    reqFork2_payload_wLen;
  reg                 _zz_reqFork1_valid;
  reg                 _zz_reqFork2_valid;
  wire                when_Stream_l945;
  wire                when_Stream_l945_1;
  wire                reqFork1_fire;
  wire                reqFork2_fire;
  wire                reqFork2_fire_1;
  wire                io_axi_w_fire;
  wire                io_axi_w_fire_1;
  reg                 cntBeat_willIncrement;
  reg                 cntBeat_willClear;
  reg        [2:0]    cntBeat_valueNext;
  reg        [2:0]    cntBeat_value;
  wire                cntBeat_willOverflowIfInc;
  wire                cntBeat_willOverflow;
  wire                io_axi_w_fire_2;
  wire                when_TxnAgent_l52;
  wire                wrDataQ_valid;
  wire                wrDataQ_ready;
  wire       [511:0]  wrDataQ_payload;
  wire                reqFork2_fire_2;
  wire                io_axi_w_fire_3;
  reg        [3:0]    _zz_wrDataQ_ready;
  wire       [1:0]    switch_Helpers_l29;
  wire                _zz_wrDataQ_ready_1;
  wire                wrDataQCtrl_valid;
  wire                wrDataQCtrl_ready;
  wire       [511:0]  wrDataQCtrl_payload;
  wire                isRdRespGrant;
  wire                when_Helpers_l40;
  wire                io_ltResp_fork2_outputs_0_valid;
  wire                io_ltResp_fork2_outputs_0_ready;
  wire       [0:0]    io_ltResp_fork2_outputs_0_payload_nId;
  wire       [21:0]   io_ltResp_fork2_outputs_0_payload_tId;
  wire       [2:0]    io_ltResp_fork2_outputs_0_payload_tabId;
  wire       [0:0]    io_ltResp_fork2_outputs_0_payload_snId;
  wire       [5:0]    io_ltResp_fork2_outputs_0_payload_txnId;
  wire       [1:0]    io_ltResp_fork2_outputs_0_payload_lkType;
  wire                io_ltResp_fork2_outputs_0_payload_lkRelease;
  wire                io_ltResp_fork2_outputs_0_payload_txnAbt;
  wire       [5:0]    io_ltResp_fork2_outputs_0_payload_lkIdx;
  wire       [2:0]    io_ltResp_fork2_outputs_0_payload_wLen;
  wire       [1:0]    io_ltResp_fork2_outputs_0_payload_respType;
  wire                io_ltResp_fork2_outputs_0_payload_lkWaited;
  wire                io_ltResp_fork2_outputs_1_valid;
  wire                io_ltResp_fork2_outputs_1_ready;
  wire       [0:0]    io_ltResp_fork2_outputs_1_payload_nId;
  wire       [21:0]   io_ltResp_fork2_outputs_1_payload_tId;
  wire       [2:0]    io_ltResp_fork2_outputs_1_payload_tabId;
  wire       [0:0]    io_ltResp_fork2_outputs_1_payload_snId;
  wire       [5:0]    io_ltResp_fork2_outputs_1_payload_txnId;
  wire       [1:0]    io_ltResp_fork2_outputs_1_payload_lkType;
  wire                io_ltResp_fork2_outputs_1_payload_lkRelease;
  wire                io_ltResp_fork2_outputs_1_payload_txnAbt;
  wire       [5:0]    io_ltResp_fork2_outputs_1_payload_lkIdx;
  wire       [2:0]    io_ltResp_fork2_outputs_1_payload_wLen;
  wire       [1:0]    io_ltResp_fork2_outputs_1_payload_respType;
  wire                io_ltResp_fork2_outputs_1_payload_lkWaited;
  reg                 _zz_io_ltResp_fork2_outputs_0_valid;
  reg                 _zz_io_ltResp_fork2_outputs_1_valid;
  wire                when_Stream_l945_2;
  wire                when_Stream_l945_3;
  wire                io_ltResp_fork2_outputs_0_fire;
  wire                io_ltResp_fork2_outputs_1_fire;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] io_ltReq_payload_lkType_string;
  reg [47:0] io_ltResp_payload_lkType_string;
  reg [71:0] io_ltResp_payload_respType_string;
  reg [47:0] lkReqQFork_payload_lkType_string;
  reg [47:0] lkReqBpss_payload_lkType_string;
  reg [47:0] _zz_io_inputs_1_payload_lkType_string;
  reg [47:0] reqFork1_payload_lkType_string;
  reg [47:0] reqFork2_payload_lkType_string;
  reg [47:0] io_ltResp_fork2_outputs_0_payload_lkType_string;
  reg [71:0] io_ltResp_fork2_outputs_0_payload_respType_string;
  reg [47:0] io_ltResp_fork2_outputs_1_payload_lkType_string;
  reg [71:0] io_ltResp_fork2_outputs_1_payload_respType_string;
  `endif


  assign _zz_io_axi_aw_payload_addr = (_zz_io_axi_aw_payload_addr_1 + 28'h0);
  assign _zz_io_axi_aw_payload_addr_1 = ({6'd0,reqFork2_payload_tId} <<< 6);
  assign _zz_io_axi_aw_payload_len = ({7'd0,1'b1} <<< reqFork2_payload_wLen);
  assign _zz_io_push_payload = (_zz_io_push_payload_1 - 8'h01);
  assign _zz_io_push_payload_1 = ({7'd0,1'b1} <<< reqFork2_payload_wLen);
  assign _zz_cntBeat_valueNext_1 = cntBeat_willIncrement;
  assign _zz_cntBeat_valueNext = {2'd0, _zz_cntBeat_valueNext_1};
  assign _zz_io_axi_ar_payload_addr = (_zz_io_axi_ar_payload_addr_1 + 28'h0);
  assign _zz_io_axi_ar_payload_addr_1 = ({6'd0,io_ltResp_payload_tId} <<< 6);
  assign _zz_io_axi_ar_payload_len = ({7'd0,1'b1} <<< io_ltResp_payload_wLen);
  StreamFifo io_lkReq_fifo (
    .io_push_valid              (io_lkReq_valid                          ), //i
    .io_push_ready              (io_lkReq_fifo_io_push_ready             ), //o
    .io_push_payload_nId        (io_lkReq_payload_nId                    ), //i
    .io_push_payload_tId        (io_lkReq_payload_tId[21:0]              ), //i
    .io_push_payload_tabId      (io_lkReq_payload_tabId[2:0]             ), //i
    .io_push_payload_snId       (io_lkReq_payload_snId                   ), //i
    .io_push_payload_txnId      (io_lkReq_payload_txnId[5:0]             ), //i
    .io_push_payload_lkType     (io_lkReq_payload_lkType[1:0]            ), //i
    .io_push_payload_lkRelease  (io_lkReq_payload_lkRelease              ), //i
    .io_push_payload_txnTimeOut (io_lkReq_payload_txnTimeOut             ), //i
    .io_push_payload_txnAbt     (io_lkReq_payload_txnAbt                 ), //i
    .io_push_payload_lkIdx      (io_lkReq_payload_lkIdx[5:0]             ), //i
    .io_push_payload_wLen       (io_lkReq_payload_wLen[2:0]              ), //i
    .io_pop_valid               (io_lkReq_fifo_io_pop_valid              ), //o
    .io_pop_ready               (streamDemux_7_io_input_ready            ), //i
    .io_pop_payload_nId         (io_lkReq_fifo_io_pop_payload_nId        ), //o
    .io_pop_payload_tId         (io_lkReq_fifo_io_pop_payload_tId[21:0]  ), //o
    .io_pop_payload_tabId       (io_lkReq_fifo_io_pop_payload_tabId[2:0] ), //o
    .io_pop_payload_snId        (io_lkReq_fifo_io_pop_payload_snId       ), //o
    .io_pop_payload_txnId       (io_lkReq_fifo_io_pop_payload_txnId[5:0] ), //o
    .io_pop_payload_lkType      (io_lkReq_fifo_io_pop_payload_lkType[1:0]), //o
    .io_pop_payload_lkRelease   (io_lkReq_fifo_io_pop_payload_lkRelease  ), //o
    .io_pop_payload_txnTimeOut  (io_lkReq_fifo_io_pop_payload_txnTimeOut ), //o
    .io_pop_payload_txnAbt      (io_lkReq_fifo_io_pop_payload_txnAbt     ), //o
    .io_pop_payload_lkIdx       (io_lkReq_fifo_io_pop_payload_lkIdx[5:0] ), //o
    .io_pop_payload_wLen        (io_lkReq_fifo_io_pop_payload_wLen[2:0]  ), //o
    .io_flush                   (1'b0                                    ), //i
    .io_occupancy               (io_lkReq_fifo_io_occupancy[3:0]         ), //o
    .io_availability            (io_lkReq_fifo_io_availability[3:0]      ), //o
    .clk                        (clk                                     ), //i
    .resetn                     (resetn                                  )  //i
  );
  StreamFifo lkReqRlseWrFifo (
    .io_push_valid              (reqFork1_valid                            ), //i
    .io_push_ready              (lkReqRlseWrFifo_io_push_ready             ), //o
    .io_push_payload_nId        (reqFork1_payload_nId                      ), //i
    .io_push_payload_tId        (reqFork1_payload_tId[21:0]                ), //i
    .io_push_payload_tabId      (reqFork1_payload_tabId[2:0]               ), //i
    .io_push_payload_snId       (reqFork1_payload_snId                     ), //i
    .io_push_payload_txnId      (reqFork1_payload_txnId[5:0]               ), //i
    .io_push_payload_lkType     (reqFork1_payload_lkType[1:0]              ), //i
    .io_push_payload_lkRelease  (reqFork1_payload_lkRelease                ), //i
    .io_push_payload_txnTimeOut (reqFork1_payload_txnTimeOut               ), //i
    .io_push_payload_txnAbt     (reqFork1_payload_txnAbt                   ), //i
    .io_push_payload_lkIdx      (reqFork1_payload_lkIdx[5:0]               ), //i
    .io_push_payload_wLen       (reqFork1_payload_wLen[2:0]                ), //i
    .io_pop_valid               (lkReqRlseWrFifo_io_pop_valid              ), //o
    .io_pop_ready               (lkReqRlseWrFifo_io_pop_ready              ), //i
    .io_pop_payload_nId         (lkReqRlseWrFifo_io_pop_payload_nId        ), //o
    .io_pop_payload_tId         (lkReqRlseWrFifo_io_pop_payload_tId[21:0]  ), //o
    .io_pop_payload_tabId       (lkReqRlseWrFifo_io_pop_payload_tabId[2:0] ), //o
    .io_pop_payload_snId        (lkReqRlseWrFifo_io_pop_payload_snId       ), //o
    .io_pop_payload_txnId       (lkReqRlseWrFifo_io_pop_payload_txnId[5:0] ), //o
    .io_pop_payload_lkType      (lkReqRlseWrFifo_io_pop_payload_lkType[1:0]), //o
    .io_pop_payload_lkRelease   (lkReqRlseWrFifo_io_pop_payload_lkRelease  ), //o
    .io_pop_payload_txnTimeOut  (lkReqRlseWrFifo_io_pop_payload_txnTimeOut ), //o
    .io_pop_payload_txnAbt      (lkReqRlseWrFifo_io_pop_payload_txnAbt     ), //o
    .io_pop_payload_lkIdx       (lkReqRlseWrFifo_io_pop_payload_lkIdx[5:0] ), //o
    .io_pop_payload_wLen        (lkReqRlseWrFifo_io_pop_payload_wLen[2:0]  ), //o
    .io_flush                   (1'b0                                      ), //i
    .io_occupancy               (lkReqRlseWrFifo_io_occupancy[3:0]         ), //o
    .io_availability            (lkReqRlseWrFifo_io_availability[3:0]      ), //o
    .clk                        (clk                                       ), //i
    .resetn                     (resetn                                    )  //i
  );
  StreamDemux streamDemux_7 (
    .io_select                       (streamDemux_7_io_select                       ), //i
    .io_input_valid                  (io_lkReq_fifo_io_pop_valid                    ), //i
    .io_input_ready                  (streamDemux_7_io_input_ready                  ), //o
    .io_input_payload_nId            (io_lkReq_fifo_io_pop_payload_nId              ), //i
    .io_input_payload_tId            (io_lkReq_fifo_io_pop_payload_tId[21:0]        ), //i
    .io_input_payload_tabId          (io_lkReq_fifo_io_pop_payload_tabId[2:0]       ), //i
    .io_input_payload_snId           (io_lkReq_fifo_io_pop_payload_snId             ), //i
    .io_input_payload_txnId          (io_lkReq_fifo_io_pop_payload_txnId[5:0]       ), //i
    .io_input_payload_lkType         (io_lkReq_fifo_io_pop_payload_lkType[1:0]      ), //i
    .io_input_payload_lkRelease      (io_lkReq_fifo_io_pop_payload_lkRelease        ), //i
    .io_input_payload_txnTimeOut     (io_lkReq_fifo_io_pop_payload_txnTimeOut       ), //i
    .io_input_payload_txnAbt         (io_lkReq_fifo_io_pop_payload_txnAbt           ), //i
    .io_input_payload_lkIdx          (io_lkReq_fifo_io_pop_payload_lkIdx[5:0]       ), //i
    .io_input_payload_wLen           (io_lkReq_fifo_io_pop_payload_wLen[2:0]        ), //i
    .io_outputs_0_valid              (streamDemux_7_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (lkReqBpss_ready                               ), //i
    .io_outputs_0_payload_nId        (streamDemux_7_io_outputs_0_payload_nId        ), //o
    .io_outputs_0_payload_tId        (streamDemux_7_io_outputs_0_payload_tId[21:0]  ), //o
    .io_outputs_0_payload_tabId      (streamDemux_7_io_outputs_0_payload_tabId[2:0] ), //o
    .io_outputs_0_payload_snId       (streamDemux_7_io_outputs_0_payload_snId       ), //o
    .io_outputs_0_payload_txnId      (streamDemux_7_io_outputs_0_payload_txnId[5:0] ), //o
    .io_outputs_0_payload_lkType     (streamDemux_7_io_outputs_0_payload_lkType[1:0]), //o
    .io_outputs_0_payload_lkRelease  (streamDemux_7_io_outputs_0_payload_lkRelease  ), //o
    .io_outputs_0_payload_txnTimeOut (streamDemux_7_io_outputs_0_payload_txnTimeOut ), //o
    .io_outputs_0_payload_txnAbt     (streamDemux_7_io_outputs_0_payload_txnAbt     ), //o
    .io_outputs_0_payload_lkIdx      (streamDemux_7_io_outputs_0_payload_lkIdx[5:0] ), //o
    .io_outputs_0_payload_wLen       (streamDemux_7_io_outputs_0_payload_wLen[2:0]  ), //o
    .io_outputs_1_valid              (streamDemux_7_io_outputs_1_valid              ), //o
    .io_outputs_1_ready              (lkReqQFork_ready                              ), //i
    .io_outputs_1_payload_nId        (streamDemux_7_io_outputs_1_payload_nId        ), //o
    .io_outputs_1_payload_tId        (streamDemux_7_io_outputs_1_payload_tId[21:0]  ), //o
    .io_outputs_1_payload_tabId      (streamDemux_7_io_outputs_1_payload_tabId[2:0] ), //o
    .io_outputs_1_payload_snId       (streamDemux_7_io_outputs_1_payload_snId       ), //o
    .io_outputs_1_payload_txnId      (streamDemux_7_io_outputs_1_payload_txnId[5:0] ), //o
    .io_outputs_1_payload_lkType     (streamDemux_7_io_outputs_1_payload_lkType[1:0]), //o
    .io_outputs_1_payload_lkRelease  (streamDemux_7_io_outputs_1_payload_lkRelease  ), //o
    .io_outputs_1_payload_txnTimeOut (streamDemux_7_io_outputs_1_payload_txnTimeOut ), //o
    .io_outputs_1_payload_txnAbt     (streamDemux_7_io_outputs_1_payload_txnAbt     ), //o
    .io_outputs_1_payload_lkIdx      (streamDemux_7_io_outputs_1_payload_lkIdx[5:0] ), //o
    .io_outputs_1_payload_wLen       (streamDemux_7_io_outputs_1_payload_wLen[2:0]  )  //o
  );
  StreamArbiter_2 streamArbiter_8 (
    .io_inputs_0_valid              (lkReqBpss_valid                              ), //i
    .io_inputs_0_ready              (streamArbiter_8_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_nId        (lkReqBpss_payload_nId                        ), //i
    .io_inputs_0_payload_tId        (lkReqBpss_payload_tId[21:0]                  ), //i
    .io_inputs_0_payload_tabId      (lkReqBpss_payload_tabId[2:0]                 ), //i
    .io_inputs_0_payload_snId       (lkReqBpss_payload_snId                       ), //i
    .io_inputs_0_payload_txnId      (lkReqBpss_payload_txnId[5:0]                 ), //i
    .io_inputs_0_payload_lkType     (lkReqBpss_payload_lkType[1:0]                ), //i
    .io_inputs_0_payload_lkRelease  (lkReqBpss_payload_lkRelease                  ), //i
    .io_inputs_0_payload_txnTimeOut (lkReqBpss_payload_txnTimeOut                 ), //i
    .io_inputs_0_payload_txnAbt     (lkReqBpss_payload_txnAbt                     ), //i
    .io_inputs_0_payload_lkIdx      (lkReqBpss_payload_lkIdx[5:0]                 ), //i
    .io_inputs_0_payload_wLen       (lkReqBpss_payload_wLen[2:0]                  ), //i
    .io_inputs_1_valid              (streamArbiter_8_io_inputs_1_valid            ), //i
    .io_inputs_1_ready              (streamArbiter_8_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_nId        (lkReqRlseWrFifo_io_pop_payload_nId           ), //i
    .io_inputs_1_payload_tId        (lkReqRlseWrFifo_io_pop_payload_tId[21:0]     ), //i
    .io_inputs_1_payload_tabId      (lkReqRlseWrFifo_io_pop_payload_tabId[2:0]    ), //i
    .io_inputs_1_payload_snId       (lkReqRlseWrFifo_io_pop_payload_snId          ), //i
    .io_inputs_1_payload_txnId      (lkReqRlseWrFifo_io_pop_payload_txnId[5:0]    ), //i
    .io_inputs_1_payload_lkType     (_zz_io_inputs_1_payload_lkType[1:0]          ), //i
    .io_inputs_1_payload_lkRelease  (lkReqRlseWrFifo_io_pop_payload_lkRelease     ), //i
    .io_inputs_1_payload_txnTimeOut (lkReqRlseWrFifo_io_pop_payload_txnTimeOut    ), //i
    .io_inputs_1_payload_txnAbt     (lkReqRlseWrFifo_io_pop_payload_txnAbt        ), //i
    .io_inputs_1_payload_lkIdx      (lkReqRlseWrFifo_io_pop_payload_lkIdx[5:0]    ), //i
    .io_inputs_1_payload_wLen       (lkReqRlseWrFifo_io_pop_payload_wLen[2:0]     ), //i
    .io_output_valid                (streamArbiter_8_io_output_valid              ), //o
    .io_output_ready                (io_ltReq_ready                               ), //i
    .io_output_payload_nId          (streamArbiter_8_io_output_payload_nId        ), //o
    .io_output_payload_tId          (streamArbiter_8_io_output_payload_tId[21:0]  ), //o
    .io_output_payload_tabId        (streamArbiter_8_io_output_payload_tabId[2:0] ), //o
    .io_output_payload_snId         (streamArbiter_8_io_output_payload_snId       ), //o
    .io_output_payload_txnId        (streamArbiter_8_io_output_payload_txnId[5:0] ), //o
    .io_output_payload_lkType       (streamArbiter_8_io_output_payload_lkType[1:0]), //o
    .io_output_payload_lkRelease    (streamArbiter_8_io_output_payload_lkRelease  ), //o
    .io_output_payload_txnTimeOut   (streamArbiter_8_io_output_payload_txnTimeOut ), //o
    .io_output_payload_txnAbt       (streamArbiter_8_io_output_payload_txnAbt     ), //o
    .io_output_payload_lkIdx        (streamArbiter_8_io_output_payload_lkIdx[5:0] ), //o
    .io_output_payload_wLen         (streamArbiter_8_io_output_payload_wLen[2:0]  ), //o
    .io_chosen                      (streamArbiter_8_io_chosen                    ), //o
    .io_chosenOH                    (streamArbiter_8_io_chosenOH[1:0]             ), //o
    .clk                            (clk                                          ), //i
    .resetn                         (resetn                                       )  //i
  );
  StreamFifoLowLatency nBeatQ (
    .io_push_valid   (reqFork2_fire_1            ), //i
    .io_push_ready   (nBeatQ_io_push_ready       ), //o
    .io_push_payload (nBeatQ_io_push_payload[2:0]), //i
    .io_pop_valid    (nBeatQ_io_pop_valid        ), //o
    .io_pop_ready    (nBeatQ_io_pop_ready        ), //i
    .io_pop_payload  (nBeatQ_io_pop_payload[2:0] ), //o
    .io_flush        (1'b0                       ), //i
    .io_occupancy    (nBeatQ_io_occupancy[3:0]   ), //o
    .clk             (clk                        ), //i
    .resetn          (resetn                     )  //i
  );
  StreamFifo_2 io_wrData_fifo (
    .io_push_valid   (io_wrData_valid                     ), //i
    .io_push_ready   (io_wrData_fifo_io_push_ready        ), //o
    .io_push_payload (io_wrData_payload[511:0]            ), //i
    .io_pop_valid    (io_wrData_fifo_io_pop_valid         ), //o
    .io_pop_ready    (wrDataQ_ready                       ), //i
    .io_pop_payload  (io_wrData_fifo_io_pop_payload[511:0]), //o
    .io_flush        (1'b0                                ), //i
    .io_occupancy    (io_wrData_fifo_io_occupancy[3:0]    ), //o
    .io_availability (io_wrData_fifo_io_availability[3:0] ), //o
    .clk             (clk                                 ), //i
    .resetn          (resetn                              )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_ltReq_payload_lkType)
      LkT_rd : io_ltReq_payload_lkType_string = "rd    ";
      LkT_wr : io_ltReq_payload_lkType_string = "wr    ";
      LkT_raw : io_ltReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_ltReq_payload_lkType_string = "insTab";
      default : io_ltReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_payload_lkType)
      LkT_rd : io_ltResp_payload_lkType_string = "rd    ";
      LkT_wr : io_ltResp_payload_lkType_string = "wr    ";
      LkT_raw : io_ltResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_ltResp_payload_lkType_string = "insTab";
      default : io_ltResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_payload_respType)
      LockRespType_grant : io_ltResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_ltResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_ltResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_ltResp_payload_respType_string = "release_1";
      default : io_ltResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(lkReqQFork_payload_lkType)
      LkT_rd : lkReqQFork_payload_lkType_string = "rd    ";
      LkT_wr : lkReqQFork_payload_lkType_string = "wr    ";
      LkT_raw : lkReqQFork_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqQFork_payload_lkType_string = "insTab";
      default : lkReqQFork_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkReqBpss_payload_lkType)
      LkT_rd : lkReqBpss_payload_lkType_string = "rd    ";
      LkT_wr : lkReqBpss_payload_lkType_string = "wr    ";
      LkT_raw : lkReqBpss_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqBpss_payload_lkType_string = "insTab";
      default : lkReqBpss_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_inputs_1_payload_lkType)
      LkT_rd : _zz_io_inputs_1_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_inputs_1_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_inputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_inputs_1_payload_lkType_string = "insTab";
      default : _zz_io_inputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(reqFork1_payload_lkType)
      LkT_rd : reqFork1_payload_lkType_string = "rd    ";
      LkT_wr : reqFork1_payload_lkType_string = "wr    ";
      LkT_raw : reqFork1_payload_lkType_string = "raw   ";
      LkT_insTab : reqFork1_payload_lkType_string = "insTab";
      default : reqFork1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(reqFork2_payload_lkType)
      LkT_rd : reqFork2_payload_lkType_string = "rd    ";
      LkT_wr : reqFork2_payload_lkType_string = "wr    ";
      LkT_raw : reqFork2_payload_lkType_string = "raw   ";
      LkT_insTab : reqFork2_payload_lkType_string = "insTab";
      default : reqFork2_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_fork2_outputs_0_payload_lkType)
      LkT_rd : io_ltResp_fork2_outputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_ltResp_fork2_outputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_ltResp_fork2_outputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_ltResp_fork2_outputs_0_payload_lkType_string = "insTab";
      default : io_ltResp_fork2_outputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_fork2_outputs_0_payload_respType)
      LockRespType_grant : io_ltResp_fork2_outputs_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_ltResp_fork2_outputs_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_ltResp_fork2_outputs_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_ltResp_fork2_outputs_0_payload_respType_string = "release_1";
      default : io_ltResp_fork2_outputs_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_fork2_outputs_1_payload_lkType)
      LkT_rd : io_ltResp_fork2_outputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_ltResp_fork2_outputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_ltResp_fork2_outputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_ltResp_fork2_outputs_1_payload_lkType_string = "insTab";
      default : io_ltResp_fork2_outputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_ltResp_fork2_outputs_1_payload_respType)
      LockRespType_grant : io_ltResp_fork2_outputs_1_payload_respType_string = "grant    ";
      LockRespType_abort : io_ltResp_fork2_outputs_1_payload_respType_string = "abort    ";
      LockRespType_waiting : io_ltResp_fork2_outputs_1_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_ltResp_fork2_outputs_1_payload_respType_string = "release_1";
      default : io_ltResp_fork2_outputs_1_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign io_lkReq_ready = io_lkReq_fifo_io_push_ready;
  assign isWrReqRlse = ((io_lkReq_fifo_io_pop_payload_lkRelease && ((io_lkReq_fifo_io_pop_payload_lkType == LkT_wr) || (io_lkReq_fifo_io_pop_payload_lkType == LkT_raw))) && (! io_lkReq_fifo_io_pop_payload_txnAbt));
  assign streamDemux_7_io_select = isWrReqRlse;
  assign lkReqBpss_valid = streamDemux_7_io_outputs_0_valid;
  assign lkReqBpss_payload_nId = streamDemux_7_io_outputs_0_payload_nId;
  assign lkReqBpss_payload_tId = streamDemux_7_io_outputs_0_payload_tId;
  assign lkReqBpss_payload_tabId = streamDemux_7_io_outputs_0_payload_tabId;
  assign lkReqBpss_payload_snId = streamDemux_7_io_outputs_0_payload_snId;
  assign lkReqBpss_payload_txnId = streamDemux_7_io_outputs_0_payload_txnId;
  assign lkReqBpss_payload_lkType = streamDemux_7_io_outputs_0_payload_lkType;
  assign lkReqBpss_payload_lkRelease = streamDemux_7_io_outputs_0_payload_lkRelease;
  assign lkReqBpss_payload_txnTimeOut = streamDemux_7_io_outputs_0_payload_txnTimeOut;
  assign lkReqBpss_payload_txnAbt = streamDemux_7_io_outputs_0_payload_txnAbt;
  assign lkReqBpss_payload_lkIdx = streamDemux_7_io_outputs_0_payload_lkIdx;
  assign lkReqBpss_payload_wLen = streamDemux_7_io_outputs_0_payload_wLen;
  assign lkReqQFork_valid = streamDemux_7_io_outputs_1_valid;
  assign lkReqQFork_payload_nId = streamDemux_7_io_outputs_1_payload_nId;
  assign lkReqQFork_payload_tId = streamDemux_7_io_outputs_1_payload_tId;
  assign lkReqQFork_payload_tabId = streamDemux_7_io_outputs_1_payload_tabId;
  assign lkReqQFork_payload_snId = streamDemux_7_io_outputs_1_payload_snId;
  assign lkReqQFork_payload_txnId = streamDemux_7_io_outputs_1_payload_txnId;
  assign lkReqQFork_payload_lkType = streamDemux_7_io_outputs_1_payload_lkType;
  assign lkReqQFork_payload_lkRelease = streamDemux_7_io_outputs_1_payload_lkRelease;
  assign lkReqQFork_payload_txnTimeOut = streamDemux_7_io_outputs_1_payload_txnTimeOut;
  assign lkReqQFork_payload_txnAbt = streamDemux_7_io_outputs_1_payload_txnAbt;
  assign lkReqQFork_payload_lkIdx = streamDemux_7_io_outputs_1_payload_lkIdx;
  assign lkReqQFork_payload_wLen = streamDemux_7_io_outputs_1_payload_wLen;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  assign lkReqRlseWrFifo_io_pop_fire = (lkReqRlseWrFifo_io_pop_valid && lkReqRlseWrFifo_io_pop_ready);
  assign switch_Helpers_l20 = {io_axi_b_fire,lkReqRlseWrFifo_io_pop_fire};
  assign _zz_io_pop_ready_1 = (4'b0000 < _zz_io_pop_ready);
  assign lkReqRlseWrFifo_io_pop_ready = (streamArbiter_8_io_inputs_1_ready && _zz_io_pop_ready_1);
  assign _zz_io_inputs_1_payload_lkType = lkReqRlseWrFifo_io_pop_payload_lkType;
  assign lkReqBpss_ready = streamArbiter_8_io_inputs_0_ready;
  assign streamArbiter_8_io_inputs_1_valid = (lkReqRlseWrFifo_io_pop_valid && _zz_io_pop_ready_1);
  assign io_ltReq_valid = streamArbiter_8_io_output_valid;
  assign io_ltReq_payload_nId = streamArbiter_8_io_output_payload_nId;
  assign io_ltReq_payload_tId = streamArbiter_8_io_output_payload_tId;
  assign io_ltReq_payload_tabId = streamArbiter_8_io_output_payload_tabId;
  assign io_ltReq_payload_snId = streamArbiter_8_io_output_payload_snId;
  assign io_ltReq_payload_txnId = streamArbiter_8_io_output_payload_txnId;
  assign io_ltReq_payload_lkType = streamArbiter_8_io_output_payload_lkType;
  assign io_ltReq_payload_lkRelease = streamArbiter_8_io_output_payload_lkRelease;
  assign io_ltReq_payload_txnTimeOut = streamArbiter_8_io_output_payload_txnTimeOut;
  assign io_ltReq_payload_txnAbt = streamArbiter_8_io_output_payload_txnAbt;
  assign io_ltReq_payload_lkIdx = streamArbiter_8_io_output_payload_lkIdx;
  assign io_ltReq_payload_wLen = streamArbiter_8_io_output_payload_wLen;
  always @(*) begin
    lkReqQFork_ready = 1'b1;
    if(when_Stream_l945) begin
      lkReqQFork_ready = 1'b0;
    end
    if(when_Stream_l945_1) begin
      lkReqQFork_ready = 1'b0;
    end
  end

  assign when_Stream_l945 = ((! reqFork1_ready) && _zz_reqFork1_valid);
  assign when_Stream_l945_1 = ((! reqFork2_ready) && _zz_reqFork2_valid);
  assign reqFork1_valid = (lkReqQFork_valid && _zz_reqFork1_valid);
  assign reqFork1_payload_nId = lkReqQFork_payload_nId;
  assign reqFork1_payload_tId = lkReqQFork_payload_tId;
  assign reqFork1_payload_tabId = lkReqQFork_payload_tabId;
  assign reqFork1_payload_snId = lkReqQFork_payload_snId;
  assign reqFork1_payload_txnId = lkReqQFork_payload_txnId;
  assign reqFork1_payload_lkType = lkReqQFork_payload_lkType;
  assign reqFork1_payload_lkRelease = lkReqQFork_payload_lkRelease;
  assign reqFork1_payload_txnTimeOut = lkReqQFork_payload_txnTimeOut;
  assign reqFork1_payload_txnAbt = lkReqQFork_payload_txnAbt;
  assign reqFork1_payload_lkIdx = lkReqQFork_payload_lkIdx;
  assign reqFork1_payload_wLen = lkReqQFork_payload_wLen;
  assign reqFork1_fire = (reqFork1_valid && reqFork1_ready);
  assign reqFork2_valid = (lkReqQFork_valid && _zz_reqFork2_valid);
  assign reqFork2_payload_nId = lkReqQFork_payload_nId;
  assign reqFork2_payload_tId = lkReqQFork_payload_tId;
  assign reqFork2_payload_tabId = lkReqQFork_payload_tabId;
  assign reqFork2_payload_snId = lkReqQFork_payload_snId;
  assign reqFork2_payload_txnId = lkReqQFork_payload_txnId;
  assign reqFork2_payload_lkType = lkReqQFork_payload_lkType;
  assign reqFork2_payload_lkRelease = lkReqQFork_payload_lkRelease;
  assign reqFork2_payload_txnTimeOut = lkReqQFork_payload_txnTimeOut;
  assign reqFork2_payload_txnAbt = lkReqQFork_payload_txnAbt;
  assign reqFork2_payload_lkIdx = lkReqQFork_payload_lkIdx;
  assign reqFork2_payload_wLen = lkReqQFork_payload_wLen;
  assign reqFork2_fire = (reqFork2_valid && reqFork2_ready);
  assign reqFork1_ready = lkReqRlseWrFifo_io_push_ready;
  assign io_axi_aw_valid = reqFork2_valid;
  assign reqFork2_ready = io_axi_aw_ready;
  assign io_axi_aw_payload_addr = {36'd0, _zz_io_axi_aw_payload_addr};
  assign io_axi_aw_payload_id = 6'h0;
  assign io_axi_aw_payload_len = (_zz_io_axi_aw_payload_len - 8'h01);
  assign io_axi_aw_payload_size = 3'b110;
  assign io_axi_aw_payload_burst = 2'b01;
  assign io_axi_w_payload_strb = 64'hffffffffffffffff;
  assign nBeatQ_io_push_payload = _zz_io_push_payload[2:0];
  assign reqFork2_fire_1 = (reqFork2_valid && reqFork2_ready);
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign nBeatQ_io_pop_ready = (io_axi_w_payload_last && io_axi_w_fire);
  assign io_axi_w_fire_1 = (io_axi_w_valid && io_axi_w_ready);
  always @(*) begin
    cntBeat_willIncrement = 1'b0;
    if(io_axi_w_fire_1) begin
      cntBeat_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    cntBeat_willClear = 1'b0;
    if(when_TxnAgent_l52) begin
      cntBeat_willClear = 1'b1;
    end
  end

  assign cntBeat_willOverflowIfInc = (cntBeat_value == 3'b111);
  assign cntBeat_willOverflow = (cntBeat_willOverflowIfInc && cntBeat_willIncrement);
  always @(*) begin
    cntBeat_valueNext = (cntBeat_value + _zz_cntBeat_valueNext);
    if(cntBeat_willClear) begin
      cntBeat_valueNext = 3'b000;
    end
  end

  assign io_axi_w_fire_2 = (io_axi_w_valid && io_axi_w_ready);
  assign when_TxnAgent_l52 = (io_axi_w_payload_last && io_axi_w_fire_2);
  assign io_wrData_ready = io_wrData_fifo_io_push_ready;
  assign wrDataQ_valid = io_wrData_fifo_io_pop_valid;
  assign wrDataQ_payload = io_wrData_fifo_io_pop_payload;
  assign reqFork2_fire_2 = (reqFork2_valid && reqFork2_ready);
  assign io_axi_w_fire_3 = (io_axi_w_valid && io_axi_w_ready);
  assign switch_Helpers_l29 = {reqFork2_fire_2,(io_axi_w_payload_last && io_axi_w_fire_3)};
  assign _zz_wrDataQ_ready_1 = (4'b0000 < _zz_wrDataQ_ready);
  assign wrDataQCtrl_valid = (wrDataQ_valid && _zz_wrDataQ_ready_1);
  assign wrDataQ_ready = (wrDataQCtrl_ready && _zz_wrDataQ_ready_1);
  assign wrDataQCtrl_payload = wrDataQ_payload;
  assign io_axi_w_payload_data = wrDataQCtrl_payload;
  assign io_axi_w_payload_last = (cntBeat_value == nBeatQ_io_pop_payload);
  assign io_axi_w_valid = wrDataQCtrl_valid;
  assign wrDataQCtrl_ready = io_axi_w_ready;
  assign io_axi_b_ready = 1'b1;
  assign isRdRespGrant = (((! io_ltResp_payload_lkRelease) && ((io_ltResp_payload_lkType == LkT_rd) || (io_ltResp_payload_lkType == LkT_raw))) && (io_ltResp_payload_respType == LockRespType_grant));
  assign when_Helpers_l40 = (! isRdRespGrant);
  always @(*) begin
    if(when_Helpers_l40) begin
      io_lkResp_valid = io_ltResp_valid;
    end else begin
      io_lkResp_valid = io_ltResp_fork2_outputs_0_valid;
    end
  end

  always @(*) begin
    if(when_Helpers_l40) begin
      io_ltResp_ready = io_lkResp_ready;
    end else begin
      io_ltResp_ready = 1'b1;
      if(when_Stream_l945_2) begin
        io_ltResp_ready = 1'b0;
      end
      if(when_Stream_l945_3) begin
        io_ltResp_ready = 1'b0;
      end
    end
  end

  always @(*) begin
    if(when_Helpers_l40) begin
      io_axi_ar_valid = 1'b0;
    end else begin
      io_axi_ar_valid = io_ltResp_fork2_outputs_1_valid;
    end
  end

  assign when_Stream_l945_2 = ((! io_ltResp_fork2_outputs_0_ready) && _zz_io_ltResp_fork2_outputs_0_valid);
  assign when_Stream_l945_3 = ((! io_ltResp_fork2_outputs_1_ready) && _zz_io_ltResp_fork2_outputs_1_valid);
  assign io_ltResp_fork2_outputs_0_valid = (io_ltResp_valid && _zz_io_ltResp_fork2_outputs_0_valid);
  assign io_ltResp_fork2_outputs_0_payload_nId = io_ltResp_payload_nId;
  assign io_ltResp_fork2_outputs_0_payload_tId = io_ltResp_payload_tId;
  assign io_ltResp_fork2_outputs_0_payload_tabId = io_ltResp_payload_tabId;
  assign io_ltResp_fork2_outputs_0_payload_snId = io_ltResp_payload_snId;
  assign io_ltResp_fork2_outputs_0_payload_txnId = io_ltResp_payload_txnId;
  assign io_ltResp_fork2_outputs_0_payload_lkType = io_ltResp_payload_lkType;
  assign io_ltResp_fork2_outputs_0_payload_lkRelease = io_ltResp_payload_lkRelease;
  assign io_ltResp_fork2_outputs_0_payload_txnAbt = io_ltResp_payload_txnAbt;
  assign io_ltResp_fork2_outputs_0_payload_lkIdx = io_ltResp_payload_lkIdx;
  assign io_ltResp_fork2_outputs_0_payload_wLen = io_ltResp_payload_wLen;
  assign io_ltResp_fork2_outputs_0_payload_respType = io_ltResp_payload_respType;
  assign io_ltResp_fork2_outputs_0_payload_lkWaited = io_ltResp_payload_lkWaited;
  assign io_ltResp_fork2_outputs_0_fire = (io_ltResp_fork2_outputs_0_valid && io_ltResp_fork2_outputs_0_ready);
  assign io_ltResp_fork2_outputs_1_valid = (io_ltResp_valid && _zz_io_ltResp_fork2_outputs_1_valid);
  assign io_ltResp_fork2_outputs_1_payload_nId = io_ltResp_payload_nId;
  assign io_ltResp_fork2_outputs_1_payload_tId = io_ltResp_payload_tId;
  assign io_ltResp_fork2_outputs_1_payload_tabId = io_ltResp_payload_tabId;
  assign io_ltResp_fork2_outputs_1_payload_snId = io_ltResp_payload_snId;
  assign io_ltResp_fork2_outputs_1_payload_txnId = io_ltResp_payload_txnId;
  assign io_ltResp_fork2_outputs_1_payload_lkType = io_ltResp_payload_lkType;
  assign io_ltResp_fork2_outputs_1_payload_lkRelease = io_ltResp_payload_lkRelease;
  assign io_ltResp_fork2_outputs_1_payload_txnAbt = io_ltResp_payload_txnAbt;
  assign io_ltResp_fork2_outputs_1_payload_lkIdx = io_ltResp_payload_lkIdx;
  assign io_ltResp_fork2_outputs_1_payload_wLen = io_ltResp_payload_wLen;
  assign io_ltResp_fork2_outputs_1_payload_respType = io_ltResp_payload_respType;
  assign io_ltResp_fork2_outputs_1_payload_lkWaited = io_ltResp_payload_lkWaited;
  assign io_ltResp_fork2_outputs_1_fire = (io_ltResp_fork2_outputs_1_valid && io_ltResp_fork2_outputs_1_ready);
  assign io_ltResp_fork2_outputs_0_ready = io_lkResp_ready;
  assign io_ltResp_fork2_outputs_1_ready = io_axi_ar_ready;
  assign io_axi_ar_payload_addr = {36'd0, _zz_io_axi_ar_payload_addr};
  assign io_axi_ar_payload_id = 6'h0;
  assign io_axi_ar_payload_len = (_zz_io_axi_ar_payload_len - 8'h01);
  assign io_axi_ar_payload_size = 3'b110;
  assign io_axi_ar_payload_burst = 2'b01;
  assign io_lkResp_payload_nId = io_ltResp_payload_nId;
  assign io_lkResp_payload_tId = io_ltResp_payload_tId;
  assign io_lkResp_payload_tabId = io_ltResp_payload_tabId;
  assign io_lkResp_payload_snId = io_ltResp_payload_snId;
  assign io_lkResp_payload_txnId = io_ltResp_payload_txnId;
  assign io_lkResp_payload_lkType = io_ltResp_payload_lkType;
  assign io_lkResp_payload_lkRelease = io_ltResp_payload_lkRelease;
  assign io_lkResp_payload_txnAbt = io_ltResp_payload_txnAbt;
  assign io_lkResp_payload_lkIdx = io_ltResp_payload_lkIdx;
  assign io_lkResp_payload_wLen = io_ltResp_payload_wLen;
  assign io_lkResp_payload_respType = io_ltResp_payload_respType;
  assign io_lkResp_payload_lkWaited = io_ltResp_payload_lkWaited;
  assign io_rdData_valid = io_axi_r_valid;
  assign io_axi_r_ready = io_rdData_ready;
  assign io_rdData_payload = io_axi_r_payload_data;
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_pop_ready <= 4'b0000;
      _zz_reqFork1_valid <= 1'b1;
      _zz_reqFork2_valid <= 1'b1;
      cntBeat_value <= 3'b000;
      _zz_wrDataQ_ready <= 4'b0000;
    end else begin
      if((switch_Helpers_l20 == {1'b1,1'b0})) begin
          _zz_io_pop_ready <= (_zz_io_pop_ready + 4'b0001);
      end else if((switch_Helpers_l20 == {1'b0,1'b1})) begin
          _zz_io_pop_ready <= (_zz_io_pop_ready - 4'b0001);
      end
      if(reqFork1_fire) begin
        _zz_reqFork1_valid <= 1'b0;
      end
      if(reqFork2_fire) begin
        _zz_reqFork2_valid <= 1'b0;
      end
      if(lkReqQFork_ready) begin
        _zz_reqFork1_valid <= 1'b1;
        _zz_reqFork2_valid <= 1'b1;
      end
      cntBeat_value <= cntBeat_valueNext;
      if((switch_Helpers_l29 == {1'b1,1'b0})) begin
          _zz_wrDataQ_ready <= (_zz_wrDataQ_ready + 4'b0001);
      end else if((switch_Helpers_l29 == {1'b0,1'b1})) begin
          _zz_wrDataQ_ready <= (_zz_wrDataQ_ready - 4'b0001);
      end
    end
  end

  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_ltResp_fork2_outputs_0_valid <= 1'b1;
      _zz_io_ltResp_fork2_outputs_1_valid <= 1'b1;
    end else begin
      if(io_ltResp_fork2_outputs_0_fire) begin
        _zz_io_ltResp_fork2_outputs_0_valid <= 1'b0;
      end
      if(io_ltResp_fork2_outputs_1_fire) begin
        _zz_io_ltResp_fork2_outputs_1_valid <= 1'b0;
      end
      if(io_ltResp_ready) begin
        _zz_io_ltResp_fork2_outputs_0_valid <= 1'b1;
        _zz_io_ltResp_fork2_outputs_1_valid <= 1'b1;
      end
    end
  end


endmodule

module LtTop (
  input      [0:0]    io_nodeId,
  input               io_lt_0_lkReq_valid,
  output              io_lt_0_lkReq_ready,
  input      [0:0]    io_lt_0_lkReq_payload_nId,
  input      [21:0]   io_lt_0_lkReq_payload_tId,
  input      [2:0]    io_lt_0_lkReq_payload_tabId,
  input      [0:0]    io_lt_0_lkReq_payload_snId,
  input      [5:0]    io_lt_0_lkReq_payload_txnId,
  input      [1:0]    io_lt_0_lkReq_payload_lkType,
  input               io_lt_0_lkReq_payload_lkRelease,
  input               io_lt_0_lkReq_payload_txnTimeOut,
  input               io_lt_0_lkReq_payload_txnAbt,
  input      [5:0]    io_lt_0_lkReq_payload_lkIdx,
  input      [2:0]    io_lt_0_lkReq_payload_wLen,
  output              io_lt_0_lkResp_valid,
  input               io_lt_0_lkResp_ready,
  output     [0:0]    io_lt_0_lkResp_payload_nId,
  output     [21:0]   io_lt_0_lkResp_payload_tId,
  output     [2:0]    io_lt_0_lkResp_payload_tabId,
  output     [0:0]    io_lt_0_lkResp_payload_snId,
  output     [5:0]    io_lt_0_lkResp_payload_txnId,
  output     [1:0]    io_lt_0_lkResp_payload_lkType,
  output              io_lt_0_lkResp_payload_lkRelease,
  output              io_lt_0_lkResp_payload_txnAbt,
  output     [5:0]    io_lt_0_lkResp_payload_lkIdx,
  output     [2:0]    io_lt_0_lkResp_payload_wLen,
  output     [1:0]    io_lt_0_lkResp_payload_respType,
  output              io_lt_0_lkResp_payload_lkWaited,
  input               io_lt_1_lkReq_valid,
  output              io_lt_1_lkReq_ready,
  input      [0:0]    io_lt_1_lkReq_payload_nId,
  input      [21:0]   io_lt_1_lkReq_payload_tId,
  input      [2:0]    io_lt_1_lkReq_payload_tabId,
  input      [0:0]    io_lt_1_lkReq_payload_snId,
  input      [5:0]    io_lt_1_lkReq_payload_txnId,
  input      [1:0]    io_lt_1_lkReq_payload_lkType,
  input               io_lt_1_lkReq_payload_lkRelease,
  input               io_lt_1_lkReq_payload_txnTimeOut,
  input               io_lt_1_lkReq_payload_txnAbt,
  input      [5:0]    io_lt_1_lkReq_payload_lkIdx,
  input      [2:0]    io_lt_1_lkReq_payload_wLen,
  output              io_lt_1_lkResp_valid,
  input               io_lt_1_lkResp_ready,
  output     [0:0]    io_lt_1_lkResp_payload_nId,
  output     [21:0]   io_lt_1_lkResp_payload_tId,
  output     [2:0]    io_lt_1_lkResp_payload_tabId,
  output     [0:0]    io_lt_1_lkResp_payload_snId,
  output     [5:0]    io_lt_1_lkResp_payload_txnId,
  output     [1:0]    io_lt_1_lkResp_payload_lkType,
  output              io_lt_1_lkResp_payload_lkRelease,
  output              io_lt_1_lkResp_payload_txnAbt,
  output     [5:0]    io_lt_1_lkResp_payload_lkIdx,
  output     [2:0]    io_lt_1_lkResp_payload_wLen,
  output     [1:0]    io_lt_1_lkResp_payload_respType,
  output              io_lt_1_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                ltChAry_0_io_lkReq_ready;
  wire                ltChAry_0_io_lkResp_valid;
  wire       [0:0]    ltChAry_0_io_lkResp_payload_nId;
  wire       [21:0]   ltChAry_0_io_lkResp_payload_tId;
  wire       [2:0]    ltChAry_0_io_lkResp_payload_tabId;
  wire       [0:0]    ltChAry_0_io_lkResp_payload_snId;
  wire       [5:0]    ltChAry_0_io_lkResp_payload_txnId;
  wire       [1:0]    ltChAry_0_io_lkResp_payload_lkType;
  wire                ltChAry_0_io_lkResp_payload_lkRelease;
  wire                ltChAry_0_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltChAry_0_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltChAry_0_io_lkResp_payload_wLen;
  wire       [1:0]    ltChAry_0_io_lkResp_payload_respType;
  wire                ltChAry_0_io_lkResp_payload_lkWaited;
  wire                streamCrossbar_2_io_inV_0_ready;
  wire                streamCrossbar_2_io_inV_1_ready;
  wire                streamCrossbar_2_io_outV_0_valid;
  wire       [0:0]    streamCrossbar_2_io_outV_0_payload_nId;
  wire       [21:0]   streamCrossbar_2_io_outV_0_payload_tId;
  wire       [2:0]    streamCrossbar_2_io_outV_0_payload_tabId;
  wire       [0:0]    streamCrossbar_2_io_outV_0_payload_snId;
  wire       [5:0]    streamCrossbar_2_io_outV_0_payload_txnId;
  wire       [1:0]    streamCrossbar_2_io_outV_0_payload_lkType;
  wire                streamCrossbar_2_io_outV_0_payload_lkRelease;
  wire                streamCrossbar_2_io_outV_0_payload_txnTimeOut;
  wire                streamCrossbar_2_io_outV_0_payload_txnAbt;
  wire       [5:0]    streamCrossbar_2_io_outV_0_payload_lkIdx;
  wire       [2:0]    streamCrossbar_2_io_outV_0_payload_wLen;
  wire                streamCrossbar_3_io_inV_0_ready;
  wire                streamCrossbar_3_io_outV_0_valid;
  wire       [0:0]    streamCrossbar_3_io_outV_0_payload_nId;
  wire       [21:0]   streamCrossbar_3_io_outV_0_payload_tId;
  wire       [2:0]    streamCrossbar_3_io_outV_0_payload_tabId;
  wire       [0:0]    streamCrossbar_3_io_outV_0_payload_snId;
  wire       [5:0]    streamCrossbar_3_io_outV_0_payload_txnId;
  wire       [1:0]    streamCrossbar_3_io_outV_0_payload_lkType;
  wire                streamCrossbar_3_io_outV_0_payload_lkRelease;
  wire                streamCrossbar_3_io_outV_0_payload_txnAbt;
  wire       [5:0]    streamCrossbar_3_io_outV_0_payload_lkIdx;
  wire       [2:0]    streamCrossbar_3_io_outV_0_payload_wLen;
  wire       [1:0]    streamCrossbar_3_io_outV_0_payload_respType;
  wire                streamCrossbar_3_io_outV_0_payload_lkWaited;
  wire                streamCrossbar_3_io_outV_1_valid;
  wire       [0:0]    streamCrossbar_3_io_outV_1_payload_nId;
  wire       [21:0]   streamCrossbar_3_io_outV_1_payload_tId;
  wire       [2:0]    streamCrossbar_3_io_outV_1_payload_tabId;
  wire       [0:0]    streamCrossbar_3_io_outV_1_payload_snId;
  wire       [5:0]    streamCrossbar_3_io_outV_1_payload_txnId;
  wire       [1:0]    streamCrossbar_3_io_outV_1_payload_lkType;
  wire                streamCrossbar_3_io_outV_1_payload_lkRelease;
  wire                streamCrossbar_3_io_outV_1_payload_txnAbt;
  wire       [5:0]    streamCrossbar_3_io_outV_1_payload_lkIdx;
  wire       [2:0]    streamCrossbar_3_io_outV_1_payload_wLen;
  wire       [1:0]    streamCrossbar_3_io_outV_1_payload_respType;
  wire                streamCrossbar_3_io_outV_1_payload_lkWaited;
  wire       [0:0]    _zz__zz_io_inDemuxSel_0;
  reg        [0:0]    _zz_io_inDemuxSel_0;
  wire                when_LtCh_l89;
  wire                when_LtCh_l92;
  `ifndef SYNTHESIS
  reg [47:0] io_lt_0_lkReq_payload_lkType_string;
  reg [47:0] io_lt_0_lkResp_payload_lkType_string;
  reg [71:0] io_lt_0_lkResp_payload_respType_string;
  reg [47:0] io_lt_1_lkReq_payload_lkType_string;
  reg [47:0] io_lt_1_lkResp_payload_lkType_string;
  reg [71:0] io_lt_1_lkResp_payload_respType_string;
  `endif


  assign _zz__zz_io_inDemuxSel_0 = (1'b1 + ltChAry_0_io_lkResp_payload_snId);
  LtCh ltChAry_0 (
    .io_lkReq_valid              (streamCrossbar_2_io_outV_0_valid              ), //i
    .io_lkReq_ready              (ltChAry_0_io_lkReq_ready                      ), //o
    .io_lkReq_payload_nId        (streamCrossbar_2_io_outV_0_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamCrossbar_2_io_outV_0_payload_tId[21:0]  ), //i
    .io_lkReq_payload_tabId      (streamCrossbar_2_io_outV_0_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamCrossbar_2_io_outV_0_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamCrossbar_2_io_outV_0_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamCrossbar_2_io_outV_0_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamCrossbar_2_io_outV_0_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamCrossbar_2_io_outV_0_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamCrossbar_2_io_outV_0_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamCrossbar_2_io_outV_0_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamCrossbar_2_io_outV_0_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltChAry_0_io_lkResp_valid                     ), //o
    .io_lkResp_ready             (streamCrossbar_3_io_inV_0_ready               ), //i
    .io_lkResp_payload_nId       (ltChAry_0_io_lkResp_payload_nId               ), //o
    .io_lkResp_payload_tId       (ltChAry_0_io_lkResp_payload_tId[21:0]         ), //o
    .io_lkResp_payload_tabId     (ltChAry_0_io_lkResp_payload_tabId[2:0]        ), //o
    .io_lkResp_payload_snId      (ltChAry_0_io_lkResp_payload_snId              ), //o
    .io_lkResp_payload_txnId     (ltChAry_0_io_lkResp_payload_txnId[5:0]        ), //o
    .io_lkResp_payload_lkType    (ltChAry_0_io_lkResp_payload_lkType[1:0]       ), //o
    .io_lkResp_payload_lkRelease (ltChAry_0_io_lkResp_payload_lkRelease         ), //o
    .io_lkResp_payload_txnAbt    (ltChAry_0_io_lkResp_payload_txnAbt            ), //o
    .io_lkResp_payload_lkIdx     (ltChAry_0_io_lkResp_payload_lkIdx[5:0]        ), //o
    .io_lkResp_payload_wLen      (ltChAry_0_io_lkResp_payload_wLen[2:0]         ), //o
    .io_lkResp_payload_respType  (ltChAry_0_io_lkResp_payload_respType[1:0]     ), //o
    .io_lkResp_payload_lkWaited  (ltChAry_0_io_lkResp_payload_lkWaited          ), //o
    .resetn                      (resetn                                        ), //i
    .clk                         (clk                                           )  //i
  );
  StreamCrossbar streamCrossbar_2 (
    .io_inV_0_valid               (io_lt_0_lkReq_valid                           ), //i
    .io_inV_0_ready               (streamCrossbar_2_io_inV_0_ready               ), //o
    .io_inV_0_payload_nId         (io_lt_0_lkReq_payload_nId                     ), //i
    .io_inV_0_payload_tId         (io_lt_0_lkReq_payload_tId[21:0]               ), //i
    .io_inV_0_payload_tabId       (io_lt_0_lkReq_payload_tabId[2:0]              ), //i
    .io_inV_0_payload_snId        (io_lt_0_lkReq_payload_snId                    ), //i
    .io_inV_0_payload_txnId       (io_lt_0_lkReq_payload_txnId[5:0]              ), //i
    .io_inV_0_payload_lkType      (io_lt_0_lkReq_payload_lkType[1:0]             ), //i
    .io_inV_0_payload_lkRelease   (io_lt_0_lkReq_payload_lkRelease               ), //i
    .io_inV_0_payload_txnTimeOut  (io_lt_0_lkReq_payload_txnTimeOut              ), //i
    .io_inV_0_payload_txnAbt      (io_lt_0_lkReq_payload_txnAbt                  ), //i
    .io_inV_0_payload_lkIdx       (io_lt_0_lkReq_payload_lkIdx[5:0]              ), //i
    .io_inV_0_payload_wLen        (io_lt_0_lkReq_payload_wLen[2:0]               ), //i
    .io_inV_1_valid               (io_lt_1_lkReq_valid                           ), //i
    .io_inV_1_ready               (streamCrossbar_2_io_inV_1_ready               ), //o
    .io_inV_1_payload_nId         (io_lt_1_lkReq_payload_nId                     ), //i
    .io_inV_1_payload_tId         (io_lt_1_lkReq_payload_tId[21:0]               ), //i
    .io_inV_1_payload_tabId       (io_lt_1_lkReq_payload_tabId[2:0]              ), //i
    .io_inV_1_payload_snId        (io_lt_1_lkReq_payload_snId                    ), //i
    .io_inV_1_payload_txnId       (io_lt_1_lkReq_payload_txnId[5:0]              ), //i
    .io_inV_1_payload_lkType      (io_lt_1_lkReq_payload_lkType[1:0]             ), //i
    .io_inV_1_payload_lkRelease   (io_lt_1_lkReq_payload_lkRelease               ), //i
    .io_inV_1_payload_txnTimeOut  (io_lt_1_lkReq_payload_txnTimeOut              ), //i
    .io_inV_1_payload_txnAbt      (io_lt_1_lkReq_payload_txnAbt                  ), //i
    .io_inV_1_payload_lkIdx       (io_lt_1_lkReq_payload_lkIdx[5:0]              ), //i
    .io_inV_1_payload_wLen        (io_lt_1_lkReq_payload_wLen[2:0]               ), //i
    .io_outV_0_valid              (streamCrossbar_2_io_outV_0_valid              ), //o
    .io_outV_0_ready              (ltChAry_0_io_lkReq_ready                      ), //i
    .io_outV_0_payload_nId        (streamCrossbar_2_io_outV_0_payload_nId        ), //o
    .io_outV_0_payload_tId        (streamCrossbar_2_io_outV_0_payload_tId[21:0]  ), //o
    .io_outV_0_payload_tabId      (streamCrossbar_2_io_outV_0_payload_tabId[2:0] ), //o
    .io_outV_0_payload_snId       (streamCrossbar_2_io_outV_0_payload_snId       ), //o
    .io_outV_0_payload_txnId      (streamCrossbar_2_io_outV_0_payload_txnId[5:0] ), //o
    .io_outV_0_payload_lkType     (streamCrossbar_2_io_outV_0_payload_lkType[1:0]), //o
    .io_outV_0_payload_lkRelease  (streamCrossbar_2_io_outV_0_payload_lkRelease  ), //o
    .io_outV_0_payload_txnTimeOut (streamCrossbar_2_io_outV_0_payload_txnTimeOut ), //o
    .io_outV_0_payload_txnAbt     (streamCrossbar_2_io_outV_0_payload_txnAbt     ), //o
    .io_outV_0_payload_lkIdx      (streamCrossbar_2_io_outV_0_payload_lkIdx[5:0] ), //o
    .io_outV_0_payload_wLen       (streamCrossbar_2_io_outV_0_payload_wLen[2:0]  ), //o
    .clk                          (clk                                           ), //i
    .resetn                       (resetn                                        )  //i
  );
  StreamCrossbar_1 streamCrossbar_3 (
    .io_inV_0_valid              (ltChAry_0_io_lkResp_valid                       ), //i
    .io_inV_0_ready              (streamCrossbar_3_io_inV_0_ready                 ), //o
    .io_inV_0_payload_nId        (ltChAry_0_io_lkResp_payload_nId                 ), //i
    .io_inV_0_payload_tId        (ltChAry_0_io_lkResp_payload_tId[21:0]           ), //i
    .io_inV_0_payload_tabId      (ltChAry_0_io_lkResp_payload_tabId[2:0]          ), //i
    .io_inV_0_payload_snId       (ltChAry_0_io_lkResp_payload_snId                ), //i
    .io_inV_0_payload_txnId      (ltChAry_0_io_lkResp_payload_txnId[5:0]          ), //i
    .io_inV_0_payload_lkType     (ltChAry_0_io_lkResp_payload_lkType[1:0]         ), //i
    .io_inV_0_payload_lkRelease  (ltChAry_0_io_lkResp_payload_lkRelease           ), //i
    .io_inV_0_payload_txnAbt     (ltChAry_0_io_lkResp_payload_txnAbt              ), //i
    .io_inV_0_payload_lkIdx      (ltChAry_0_io_lkResp_payload_lkIdx[5:0]          ), //i
    .io_inV_0_payload_wLen       (ltChAry_0_io_lkResp_payload_wLen[2:0]           ), //i
    .io_inV_0_payload_respType   (ltChAry_0_io_lkResp_payload_respType[1:0]       ), //i
    .io_inV_0_payload_lkWaited   (ltChAry_0_io_lkResp_payload_lkWaited            ), //i
    .io_outV_0_valid             (streamCrossbar_3_io_outV_0_valid                ), //o
    .io_outV_0_ready             (io_lt_0_lkResp_ready                            ), //i
    .io_outV_0_payload_nId       (streamCrossbar_3_io_outV_0_payload_nId          ), //o
    .io_outV_0_payload_tId       (streamCrossbar_3_io_outV_0_payload_tId[21:0]    ), //o
    .io_outV_0_payload_tabId     (streamCrossbar_3_io_outV_0_payload_tabId[2:0]   ), //o
    .io_outV_0_payload_snId      (streamCrossbar_3_io_outV_0_payload_snId         ), //o
    .io_outV_0_payload_txnId     (streamCrossbar_3_io_outV_0_payload_txnId[5:0]   ), //o
    .io_outV_0_payload_lkType    (streamCrossbar_3_io_outV_0_payload_lkType[1:0]  ), //o
    .io_outV_0_payload_lkRelease (streamCrossbar_3_io_outV_0_payload_lkRelease    ), //o
    .io_outV_0_payload_txnAbt    (streamCrossbar_3_io_outV_0_payload_txnAbt       ), //o
    .io_outV_0_payload_lkIdx     (streamCrossbar_3_io_outV_0_payload_lkIdx[5:0]   ), //o
    .io_outV_0_payload_wLen      (streamCrossbar_3_io_outV_0_payload_wLen[2:0]    ), //o
    .io_outV_0_payload_respType  (streamCrossbar_3_io_outV_0_payload_respType[1:0]), //o
    .io_outV_0_payload_lkWaited  (streamCrossbar_3_io_outV_0_payload_lkWaited     ), //o
    .io_outV_1_valid             (streamCrossbar_3_io_outV_1_valid                ), //o
    .io_outV_1_ready             (io_lt_1_lkResp_ready                            ), //i
    .io_outV_1_payload_nId       (streamCrossbar_3_io_outV_1_payload_nId          ), //o
    .io_outV_1_payload_tId       (streamCrossbar_3_io_outV_1_payload_tId[21:0]    ), //o
    .io_outV_1_payload_tabId     (streamCrossbar_3_io_outV_1_payload_tabId[2:0]   ), //o
    .io_outV_1_payload_snId      (streamCrossbar_3_io_outV_1_payload_snId         ), //o
    .io_outV_1_payload_txnId     (streamCrossbar_3_io_outV_1_payload_txnId[5:0]   ), //o
    .io_outV_1_payload_lkType    (streamCrossbar_3_io_outV_1_payload_lkType[1:0]  ), //o
    .io_outV_1_payload_lkRelease (streamCrossbar_3_io_outV_1_payload_lkRelease    ), //o
    .io_outV_1_payload_txnAbt    (streamCrossbar_3_io_outV_1_payload_txnAbt       ), //o
    .io_outV_1_payload_lkIdx     (streamCrossbar_3_io_outV_1_payload_lkIdx[5:0]   ), //o
    .io_outV_1_payload_wLen      (streamCrossbar_3_io_outV_1_payload_wLen[2:0]    ), //o
    .io_outV_1_payload_respType  (streamCrossbar_3_io_outV_1_payload_respType[1:0]), //o
    .io_outV_1_payload_lkWaited  (streamCrossbar_3_io_outV_1_payload_lkWaited     ), //o
    .io_inDemuxSel_0             (_zz_io_inDemuxSel_0                             ), //i
    .clk                         (clk                                             ), //i
    .resetn                      (resetn                                          )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lt_0_lkReq_payload_lkType)
      LkT_rd : io_lt_0_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lt_0_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lt_0_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lt_0_lkReq_payload_lkType_string = "insTab";
      default : io_lt_0_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lt_0_lkResp_payload_lkType)
      LkT_rd : io_lt_0_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lt_0_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lt_0_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lt_0_lkResp_payload_lkType_string = "insTab";
      default : io_lt_0_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lt_0_lkResp_payload_respType)
      LockRespType_grant : io_lt_0_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lt_0_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lt_0_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lt_0_lkResp_payload_respType_string = "release_1";
      default : io_lt_0_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_lt_1_lkReq_payload_lkType)
      LkT_rd : io_lt_1_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lt_1_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lt_1_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lt_1_lkReq_payload_lkType_string = "insTab";
      default : io_lt_1_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lt_1_lkResp_payload_lkType)
      LkT_rd : io_lt_1_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lt_1_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lt_1_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lt_1_lkResp_payload_lkType_string = "insTab";
      default : io_lt_1_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lt_1_lkResp_payload_respType)
      LockRespType_grant : io_lt_1_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lt_1_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lt_1_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lt_1_lkResp_payload_respType_string = "release_1";
      default : io_lt_1_lkResp_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign io_lt_0_lkReq_ready = streamCrossbar_2_io_inV_0_ready;
  assign io_lt_1_lkReq_ready = streamCrossbar_2_io_inV_1_ready;
  assign when_LtCh_l89 = (io_nodeId < ltChAry_0_io_lkResp_payload_snId);
  always @(*) begin
    if(when_LtCh_l89) begin
      _zz_io_inDemuxSel_0 = (_zz__zz_io_inDemuxSel_0 - 1'b1);
    end else begin
      if(when_LtCh_l92) begin
        _zz_io_inDemuxSel_0 = (1'b1 + ltChAry_0_io_lkResp_payload_snId);
      end else begin
        _zz_io_inDemuxSel_0 = 1'b0;
      end
    end
  end

  assign when_LtCh_l92 = (ltChAry_0_io_lkResp_payload_snId < io_nodeId);
  assign io_lt_0_lkResp_valid = streamCrossbar_3_io_outV_0_valid;
  assign io_lt_0_lkResp_payload_nId = streamCrossbar_3_io_outV_0_payload_nId;
  assign io_lt_0_lkResp_payload_tId = streamCrossbar_3_io_outV_0_payload_tId;
  assign io_lt_0_lkResp_payload_tabId = streamCrossbar_3_io_outV_0_payload_tabId;
  assign io_lt_0_lkResp_payload_snId = streamCrossbar_3_io_outV_0_payload_snId;
  assign io_lt_0_lkResp_payload_txnId = streamCrossbar_3_io_outV_0_payload_txnId;
  assign io_lt_0_lkResp_payload_lkType = streamCrossbar_3_io_outV_0_payload_lkType;
  assign io_lt_0_lkResp_payload_lkRelease = streamCrossbar_3_io_outV_0_payload_lkRelease;
  assign io_lt_0_lkResp_payload_txnAbt = streamCrossbar_3_io_outV_0_payload_txnAbt;
  assign io_lt_0_lkResp_payload_lkIdx = streamCrossbar_3_io_outV_0_payload_lkIdx;
  assign io_lt_0_lkResp_payload_wLen = streamCrossbar_3_io_outV_0_payload_wLen;
  assign io_lt_0_lkResp_payload_respType = streamCrossbar_3_io_outV_0_payload_respType;
  assign io_lt_0_lkResp_payload_lkWaited = streamCrossbar_3_io_outV_0_payload_lkWaited;
  assign io_lt_1_lkResp_valid = streamCrossbar_3_io_outV_1_valid;
  assign io_lt_1_lkResp_payload_nId = streamCrossbar_3_io_outV_1_payload_nId;
  assign io_lt_1_lkResp_payload_tId = streamCrossbar_3_io_outV_1_payload_tId;
  assign io_lt_1_lkResp_payload_tabId = streamCrossbar_3_io_outV_1_payload_tabId;
  assign io_lt_1_lkResp_payload_snId = streamCrossbar_3_io_outV_1_payload_snId;
  assign io_lt_1_lkResp_payload_txnId = streamCrossbar_3_io_outV_1_payload_txnId;
  assign io_lt_1_lkResp_payload_lkType = streamCrossbar_3_io_outV_1_payload_lkType;
  assign io_lt_1_lkResp_payload_lkRelease = streamCrossbar_3_io_outV_1_payload_lkRelease;
  assign io_lt_1_lkResp_payload_txnAbt = streamCrossbar_3_io_outV_1_payload_txnAbt;
  assign io_lt_1_lkResp_payload_lkIdx = streamCrossbar_3_io_outV_1_payload_lkIdx;
  assign io_lt_1_lkResp_payload_wLen = streamCrossbar_3_io_outV_1_payload_wLen;
  assign io_lt_1_lkResp_payload_respType = streamCrossbar_3_io_outV_1_payload_respType;
  assign io_lt_1_lkResp_payload_lkWaited = streamCrossbar_3_io_outV_1_payload_lkWaited;

endmodule

module TxnManCS (
  output              io_lkReqLoc_valid,
  input               io_lkReqLoc_ready,
  output     [0:0]    io_lkReqLoc_payload_nId,
  output     [21:0]   io_lkReqLoc_payload_tId,
  output     [2:0]    io_lkReqLoc_payload_tabId,
  output     [0:0]    io_lkReqLoc_payload_snId,
  output     [5:0]    io_lkReqLoc_payload_txnId,
  output     [1:0]    io_lkReqLoc_payload_lkType,
  output              io_lkReqLoc_payload_lkRelease,
  output              io_lkReqLoc_payload_txnTimeOut,
  output              io_lkReqLoc_payload_txnAbt,
  output     [5:0]    io_lkReqLoc_payload_lkIdx,
  output     [2:0]    io_lkReqLoc_payload_wLen,
  output              io_lkReqRmt_valid,
  input               io_lkReqRmt_ready,
  output     [0:0]    io_lkReqRmt_payload_nId,
  output     [21:0]   io_lkReqRmt_payload_tId,
  output     [2:0]    io_lkReqRmt_payload_tabId,
  output     [0:0]    io_lkReqRmt_payload_snId,
  output     [5:0]    io_lkReqRmt_payload_txnId,
  output     [1:0]    io_lkReqRmt_payload_lkType,
  output              io_lkReqRmt_payload_lkRelease,
  output              io_lkReqRmt_payload_txnTimeOut,
  output              io_lkReqRmt_payload_txnAbt,
  output     [5:0]    io_lkReqRmt_payload_lkIdx,
  output     [2:0]    io_lkReqRmt_payload_wLen,
  input               io_lkRespLoc_valid,
  output              io_lkRespLoc_ready,
  input      [0:0]    io_lkRespLoc_payload_nId,
  input      [21:0]   io_lkRespLoc_payload_tId,
  input      [2:0]    io_lkRespLoc_payload_tabId,
  input      [0:0]    io_lkRespLoc_payload_snId,
  input      [5:0]    io_lkRespLoc_payload_txnId,
  input      [1:0]    io_lkRespLoc_payload_lkType,
  input               io_lkRespLoc_payload_lkRelease,
  input               io_lkRespLoc_payload_txnAbt,
  input      [5:0]    io_lkRespLoc_payload_lkIdx,
  input      [2:0]    io_lkRespLoc_payload_wLen,
  input      [1:0]    io_lkRespLoc_payload_respType,
  input               io_lkRespLoc_payload_lkWaited,
  input               io_lkRespRmt_valid,
  output              io_lkRespRmt_ready,
  input      [0:0]    io_lkRespRmt_payload_nId,
  input      [21:0]   io_lkRespRmt_payload_tId,
  input      [2:0]    io_lkRespRmt_payload_tabId,
  input      [0:0]    io_lkRespRmt_payload_snId,
  input      [5:0]    io_lkRespRmt_payload_txnId,
  input      [1:0]    io_lkRespRmt_payload_lkType,
  input               io_lkRespRmt_payload_lkRelease,
  input               io_lkRespRmt_payload_txnAbt,
  input      [5:0]    io_lkRespRmt_payload_lkIdx,
  input      [2:0]    io_lkRespRmt_payload_wLen,
  input      [1:0]    io_lkRespRmt_payload_respType,
  input               io_lkRespRmt_payload_lkWaited,
  input               io_rdRmt_valid,
  output              io_rdRmt_ready,
  input      [511:0]  io_rdRmt_payload,
  output              io_wrRmt_valid,
  input               io_wrRmt_ready,
  output     [511:0]  io_wrRmt_payload,
  output              io_axi_aw_valid,
  input               io_axi_aw_ready,
  output     [63:0]   io_axi_aw_payload_addr,
  output     [5:0]    io_axi_aw_payload_id,
  output     [7:0]    io_axi_aw_payload_len,
  output     [2:0]    io_axi_aw_payload_size,
  output     [1:0]    io_axi_aw_payload_burst,
  output              io_axi_w_valid,
  input               io_axi_w_ready,
  output     [511:0]  io_axi_w_payload_data,
  output     [63:0]   io_axi_w_payload_strb,
  output              io_axi_w_payload_last,
  input               io_axi_b_valid,
  output              io_axi_b_ready,
  input      [5:0]    io_axi_b_payload_id,
  input      [1:0]    io_axi_b_payload_resp,
  output              io_axi_ar_valid,
  input               io_axi_ar_ready,
  output     [63:0]   io_axi_ar_payload_addr,
  output     [5:0]    io_axi_ar_payload_id,
  output     [7:0]    io_axi_ar_payload_len,
  output     [2:0]    io_axi_ar_payload_size,
  output     [1:0]    io_axi_ar_payload_burst,
  input               io_axi_r_valid,
  output              io_axi_r_ready,
  input      [511:0]  io_axi_r_payload_data,
  input      [5:0]    io_axi_r_payload_id,
  input      [1:0]    io_axi_r_payload_resp,
  input               io_axi_r_payload_last,
  output              io_cmdAxi_aw_valid,
  input               io_cmdAxi_aw_ready,
  output     [63:0]   io_cmdAxi_aw_payload_addr,
  output     [5:0]    io_cmdAxi_aw_payload_id,
  output     [7:0]    io_cmdAxi_aw_payload_len,
  output     [2:0]    io_cmdAxi_aw_payload_size,
  output     [1:0]    io_cmdAxi_aw_payload_burst,
  output              io_cmdAxi_w_valid,
  input               io_cmdAxi_w_ready,
  output     [511:0]  io_cmdAxi_w_payload_data,
  output     [63:0]   io_cmdAxi_w_payload_strb,
  output              io_cmdAxi_w_payload_last,
  input               io_cmdAxi_b_valid,
  output              io_cmdAxi_b_ready,
  input      [5:0]    io_cmdAxi_b_payload_id,
  input      [1:0]    io_cmdAxi_b_payload_resp,
  output              io_cmdAxi_ar_valid,
  input               io_cmdAxi_ar_ready,
  output     [63:0]   io_cmdAxi_ar_payload_addr,
  output     [5:0]    io_cmdAxi_ar_payload_id,
  output     [7:0]    io_cmdAxi_ar_payload_len,
  output     [2:0]    io_cmdAxi_ar_payload_size,
  output     [1:0]    io_cmdAxi_ar_payload_burst,
  input               io_cmdAxi_r_valid,
  output              io_cmdAxi_r_ready,
  input      [511:0]  io_cmdAxi_r_payload_data,
  input      [5:0]    io_cmdAxi_r_payload_id,
  input      [1:0]    io_cmdAxi_r_payload_resp,
  input               io_cmdAxi_r_payload_last,
  input               io_start,
  input      [0:0]    io_nodeId,
  input      [31:0]   io_txnNumTotal,
  input      [31:0]   io_cmdAddrOffs,
  output reg          io_done,
  output reg [31:0]   io_cntTxnCmt,
  output reg [31:0]   io_cntTxnAbt,
  output reg [31:0]   io_cntTxnLd,
  output reg [31:0]   io_cntLockLoc,
  output reg [31:0]   io_cntLockRmt,
  output reg [31:0]   io_cntLockDenyLoc,
  output reg [31:0]   io_cntLockDenyRmt,
  output reg [31:0]   io_cntClk,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam compLkRespLoc_enumDef_BOOT = 2'd0;
  localparam compLkRespLoc_enumDef_WAIT_RESP = 2'd1;
  localparam compLkRespLoc_enumDef_LOCAL_RD_REQ = 2'd2;
  localparam compLkRespRmt_enumDef_BOOT = 2'd0;
  localparam compLkRespRmt_enumDef_WAIT_RESP = 2'd1;
  localparam compLkRespRmt_enumDef_RMT_RD_CONSUME = 2'd2;
  localparam compTxnCmtLoc_enumDef_BOOT = 2'd0;
  localparam compTxnCmtLoc_enumDef_CS_TXN = 2'd1;
  localparam compTxnCmtLoc_enumDef_LOCAL_AW = 2'd2;
  localparam compTxnCmtLoc_enumDef_LOCAL_W = 2'd3;
  localparam compLkRlseRmt_enumDef_BOOT = 2'd0;
  localparam compLkRlseRmt_enumDef_CS_TXN = 2'd1;
  localparam compLkRlseRmt_enumDef_RMT_LK_RLSE = 2'd2;
  localparam compLkRlseRmt_enumDef_RMT_WR = 2'd3;
  localparam compLoadTxn_enumDef_BOOT = 3'd0;
  localparam compLoadTxn_enumDef_IDLE = 3'd1;
  localparam compLoadTxn_enumDef_CS_TXN = 3'd2;
  localparam compLoadTxn_enumDef_RD_CMDAXI = 3'd3;
  localparam compLoadTxn_enumDef_LD_TXN = 3'd4;
  localparam compLkReq_enumDef_BOOT = 2'd0;
  localparam compLkReq_enumDef_CS_TXN = 2'd1;
  localparam compLkReq_enumDef_RD_TXN = 2'd2;
  localparam compLkRlseLoc_enumDef_BOOT = 2'd0;
  localparam compLkRlseLoc_enumDef_CS_TXN = 2'd1;
  localparam compLkRlseLoc_enumDef_LK_RLSE = 2'd2;
  localparam compTimeOut_enumDef_BOOT = 2'd0;
  localparam compTimeOut_enumDef_IDLE = 2'd1;
  localparam compTimeOut_enumDef_COUNT = 2'd2;
  localparam clkCnt_enumDef_BOOT = 2'd0;
  localparam clkCnt_enumDef_IDLE = 2'd1;
  localparam clkCnt_enumDef_CNT = 2'd2;

  wire                streamArbiter_8_io_output_ready;
  wire                streamArbiter_9_io_output_ready;
  reg        [30:0]   _zz_txnMem_port0;
  reg        [30:0]   _zz_txnWrMemLoc_port0;
  reg        [48:0]   _zz_lkMemLoc_port0;
  reg        [48:0]   _zz_lkMemRmt_port0;
  wire                streamArbiter_8_io_inputs_0_ready;
  wire                streamArbiter_8_io_inputs_1_ready;
  wire                streamArbiter_8_io_output_valid;
  wire       [0:0]    streamArbiter_8_io_output_payload_nId;
  wire       [21:0]   streamArbiter_8_io_output_payload_tId;
  wire       [2:0]    streamArbiter_8_io_output_payload_tabId;
  wire       [0:0]    streamArbiter_8_io_output_payload_snId;
  wire       [5:0]    streamArbiter_8_io_output_payload_txnId;
  wire       [1:0]    streamArbiter_8_io_output_payload_lkType;
  wire                streamArbiter_8_io_output_payload_lkRelease;
  wire                streamArbiter_8_io_output_payload_txnTimeOut;
  wire                streamArbiter_8_io_output_payload_txnAbt;
  wire       [5:0]    streamArbiter_8_io_output_payload_lkIdx;
  wire       [2:0]    streamArbiter_8_io_output_payload_wLen;
  wire       [0:0]    streamArbiter_8_io_chosen;
  wire       [1:0]    streamArbiter_8_io_chosenOH;
  wire                streamArbiter_9_io_inputs_0_ready;
  wire                streamArbiter_9_io_inputs_1_ready;
  wire                streamArbiter_9_io_output_valid;
  wire       [0:0]    streamArbiter_9_io_output_payload_nId;
  wire       [21:0]   streamArbiter_9_io_output_payload_tId;
  wire       [2:0]    streamArbiter_9_io_output_payload_tabId;
  wire       [0:0]    streamArbiter_9_io_output_payload_snId;
  wire       [5:0]    streamArbiter_9_io_output_payload_txnId;
  wire       [1:0]    streamArbiter_9_io_output_payload_lkType;
  wire                streamArbiter_9_io_output_payload_lkRelease;
  wire                streamArbiter_9_io_output_payload_txnTimeOut;
  wire                streamArbiter_9_io_output_payload_txnAbt;
  wire       [5:0]    streamArbiter_9_io_output_payload_lkIdx;
  wire       [2:0]    streamArbiter_9_io_output_payload_wLen;
  wire       [0:0]    streamArbiter_9_io_chosen;
  wire       [1:0]    streamArbiter_9_io_chosenOH;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start;
  wire       [58:0]   _zz_compLkReq_mskTxn2Start_1;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_2;
  wire       [52:0]   _zz_compLkReq_mskTxn2Start_3;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_4;
  wire       [46:0]   _zz_compLkReq_mskTxn2Start_5;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_6;
  wire       [40:0]   _zz_compLkReq_mskTxn2Start_7;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_8;
  wire       [34:0]   _zz_compLkReq_mskTxn2Start_9;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_10;
  wire       [28:0]   _zz_compLkReq_mskTxn2Start_11;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_12;
  wire       [22:0]   _zz_compLkReq_mskTxn2Start_13;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_14;
  wire       [16:0]   _zz_compLkReq_mskTxn2Start_15;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_16;
  wire       [10:0]   _zz_compLkReq_mskTxn2Start_17;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_18;
  wire       [4:0]    _zz_compLkReq_mskTxn2Start_19;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_20;
  wire       [58:0]   _zz_compLkReq_mskTxn2Start_21;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_22;
  wire       [52:0]   _zz_compLkReq_mskTxn2Start_23;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_24;
  wire       [46:0]   _zz_compLkReq_mskTxn2Start_25;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_26;
  wire       [40:0]   _zz_compLkReq_mskTxn2Start_27;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_28;
  wire       [34:0]   _zz_compLkReq_mskTxn2Start_29;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_30;
  wire       [28:0]   _zz_compLkReq_mskTxn2Start_31;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_32;
  wire       [22:0]   _zz_compLkReq_mskTxn2Start_33;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_34;
  wire       [16:0]   _zz_compLkReq_mskTxn2Start_35;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_36;
  wire       [10:0]   _zz_compLkReq_mskTxn2Start_37;
  wire       [0:0]    _zz_compLkReq_mskTxn2Start_38;
  wire       [4:0]    _zz_compLkReq_mskTxn2Start_39;
  wire       [63:0]   _zz_compLkReq_mskTxn2Start_ohFirst_masked;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_57;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_58;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_59;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_60;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_61;
  wire                _zz__zz_compLkReq_rIdxTxn2Start_62;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlse;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlse_1;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlse_2;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlse_3;
  reg        [5:0]    _zz_compLkRespLoc_getAllLkResp;
  reg        [5:0]    _zz_compLkRespLoc_getAllLkResp_1;
  reg        [5:0]    _zz_compLkRespLoc_getAllLkResp_2;
  reg        [5:0]    _zz_compLkRespLoc_getAllLkResp_3;
  reg        [5:0]    _zz__zz_cntRlseRespLoc_0;
  reg        [5:0]    _zz__zz_cntLkHoldLoc_0;
  reg        [5:0]    _zz__zz_cntLkWaitLoc_0;
  wire       [5:0]    _zz_compLkRespLoc_getAllRlseTimeOut;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlseTimeOut_1;
  wire       [5:0]    _zz_compLkRespLoc_getAllRlseTimeOut_2;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlseTimeOut_3;
  reg        [5:0]    _zz_compLkRespLoc_getAllRlseTimeOut_4;
  reg                 _zz_when_TxnManCS_l166;
  reg                 _zz_when_TxnManCS_l164;
  reg                 _zz_when_TxnManCS_l164_1;
  wire       [27:0]   _zz_io_axi_ar_payload_addr;
  wire       [27:0]   _zz_io_axi_ar_payload_addr_1;
  wire       [7:0]    _zz_io_axi_ar_payload_len;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlse;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlse_1;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlse_2;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlse_3;
  reg        [5:0]    _zz_compLkRespRmt_getAllLkResp;
  reg        [5:0]    _zz_compLkRespRmt_getAllLkResp_1;
  reg        [5:0]    _zz_compLkRespRmt_getAllLkResp_2;
  reg        [5:0]    _zz_compLkRespRmt_getAllLkResp_3;
  reg        [5:0]    _zz__zz_cntRlseRespRmt_0;
  reg        [5:0]    _zz__zz_cntLkHoldRmt_0;
  reg        [5:0]    _zz__zz_cntLkWaitRmt_0;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlseTimeOut;
  wire       [5:0]    _zz_compLkRespRmt_getAllRlseTimeOut_1;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlseTimeOut_2;
  reg        [5:0]    _zz_compLkRespRmt_getAllRlseTimeOut_3;
  wire       [5:0]    _zz_compLkRespRmt_getAllRlseTimeOut_4;
  reg                 _zz_when_TxnManCS_l261;
  reg                 _zz_when_TxnManCS_l259;
  reg                 _zz_when_TxnManCS_l259_1;
  reg        [5:0]    _zz__zz_cntCmtRespLoc_0;
  reg        [5:0]    _zz__zz_cntCmtReqLoc_0;
  wire       [11:0]   _zz__zz_compTxnCmtLoc_cmtTxn_nId;
  wire                _zz_txnWrMemLoc_port;
  wire                _zz__zz_compTxnCmtLoc_cmtTxn_nId_1;
  reg        [5:0]    _zz_compTxnCmtLoc_getAllLkResp;
  reg        [5:0]    _zz_compTxnCmtLoc_getAllLkResp_1;
  reg        [5:0]    _zz_compTxnCmtLoc_getAllLkResp_2;
  reg        [5:0]    _zz_compTxnCmtLoc_getAllLkResp_3;
  wire       [27:0]   _zz_io_axi_aw_payload_addr;
  wire       [27:0]   _zz_io_axi_aw_payload_addr_1;
  wire       [7:0]    _zz_io_axi_aw_payload_len;
  wire       [7:0]    _zz_io_axi_w_payload_last;
  wire       [7:0]    _zz_io_axi_w_payload_last_1;
  reg        [5:0]    _zz__zz_cntRlseReqLoc_0;
  wire       [11:0]   _zz__zz_compLkRlseLoc_lkItem_nId;
  wire                _zz_lkMemLoc_port;
  wire                _zz__zz_compLkRlseLoc_lkItem_nId_1;
  reg        [5:0]    _zz_compLkRlseLoc_getAllLkResp;
  reg        [5:0]    _zz_compLkRlseLoc_getAllLkResp_1;
  reg        [5:0]    _zz_compLkRlseLoc_getAllLkResp_2;
  reg        [5:0]    _zz_compLkRlseLoc_getAllLkResp_3;
  reg                 _zz__zz_lkReqRlseLoc_payload_txnAbt;
  reg                 _zz__zz_lkReqRlseLoc_payload_txnTimeOut;
  reg        [5:0]    _zz__zz_cntRlseReqRmt_0;
  wire       [11:0]   _zz__zz_compLkRlseRmt_lkItem_nId;
  wire                _zz_lkMemRmt_port;
  wire                _zz__zz_compLkRlseRmt_lkItem_nId_1;
  reg        [5:0]    _zz_compLkRlseRmt_getAllLkResp;
  reg        [5:0]    _zz_compLkRlseRmt_getAllLkResp_1;
  reg        [5:0]    _zz_compLkRlseRmt_getAllLkResp_2;
  reg        [5:0]    _zz_compLkRlseRmt_getAllLkResp_3;
  reg                 _zz__zz_lkReqRlseRmt_payload_txnAbt;
  reg                 _zz__zz_lkReqRlseRmt_payload_txnTimeOut;
  wire       [40:0]   _zz_io_cmdAxi_ar_payload_addr;
  wire       [40:0]   _zz_io_cmdAxi_ar_payload_addr_1;
  wire       [37:0]   _zz_io_cmdAxi_ar_payload_addr_2;
  wire       [40:0]   _zz_io_cmdAxi_ar_payload_addr_3;
  wire       [37:0]   _zz_io_cmdAxi_ar_payload_addr_4;
  wire       [3:0]    _zz_io_cmdAxi_ar_payload_len;
  wire       [3:0]    _zz_io_cmdAxi_ar_payload_len_1;
  wire       [2:0]    _zz_compLoadTxn_cntTxnWordInLine_valueNext;
  wire       [0:0]    _zz_compLoadTxn_cntTxnWordInLine_valueNext_1;
  wire       [5:0]    _zz_compLoadTxn_cntTxnWord_valueNext;
  wire       [0:0]    _zz_compLoadTxn_cntTxnWord_valueNext_1;
  reg        [63:0]   _zz_compLoadTxn_bitsBuff;
  wire                _zz_when_TxnManCS_l672;
  wire                _zz_when_TxnManCS_l672_1;
  wire                _zz_when_TxnManCS_l672_2;
  wire                _zz_when_TxnManCS_l672_3;
  wire       [11:0]   _zz_txnWrMemLoc_port_1;
  wire       [11:0]   _zz_txnWrMemLoc_port_2;
  wire       [30:0]   _zz_txnWrMemLoc_port_3;
  wire       [11:0]   _zz_txnWrMemRmt_port;
  wire       [11:0]   _zz_txnWrMemRmt_port_1;
  wire       [30:0]   _zz_txnWrMemRmt_port_2;
  wire       [30:0]   _zz_compLkReq_txnLen;
  wire       [11:0]   _zz__zz_compLkReq_txnMemRdCmd_payload;
  wire       [11:0]   _zz__zz_compLkReq_txnMemRdCmd_payload_1;
  wire       [11:0]   _zz_compLkReq_txnMemRdCmd_payload_1;
  reg        [5:0]    _zz__zz_cntLkReqLoc_0;
  reg        [5:0]    _zz__zz_cntLkReqRmt_0;
  reg        [5:0]    _zz__zz_cntLkReqWrLoc_0;
  reg        [5:0]    _zz__zz_cntLkReqWrRmt_0;
  wire       [5:0]    _zz_when_TxnManCS_l128;
  reg                 _zz_when_TxnManCS_l128_1;
  wire       [11:0]   _zz_lkMemLoc_port_1;
  wire       [11:0]   _zz_lkMemLoc_port_2;
  wire       [11:0]   _zz_lkMemLoc_port_3;
  wire       [11:0]   _zz_lkMemLoc_port_4;
  wire       [48:0]   _zz_lkMemLoc_port_5;
  reg        [5:0]    _zz__zz_cntLkRespLoc_0;
  reg        [5:0]    _zz__zz_cntLkHoldWrLoc_0;
  wire       [11:0]   _zz_lkMemRmt_port_1;
  wire       [11:0]   _zz_lkMemRmt_port_2;
  wire       [11:0]   _zz_lkMemRmt_port_3;
  wire       [11:0]   _zz_lkMemRmt_port_4;
  wire       [48:0]   _zz_lkMemRmt_port_5;
  reg        [5:0]    _zz__zz_cntLkRespRmt_0;
  reg        [5:0]    _zz__zz_cntLkHoldWrRmt_0;
  wire       [7:0]    _zz_when_TxnManCS_l315;
  wire       [7:0]    _zz_when_TxnManCS_l315_1;
  reg                 _zz_when_TxnManCS_l369;
  reg                 _zz_when_TxnManCS_l369_1;
  reg        [5:0]    _zz_when_TxnManCS_l369_2;
  reg        [5:0]    _zz__zz_cntRlseReqWrLoc_0;
  reg        [5:0]    _zz__zz_when_TxnManCS_l440;
  reg                 _zz_when_TxnManCS_l440_1;
  reg        [5:0]    _zz_when_TxnManCS_l440_2;
  wire       [5:0]    _zz_when_TxnManCS_l440_3;
  reg        [5:0]    _zz_when_TxnManCS_l440_4;
  reg        [5:0]    _zz__zz_when_TxnManCS_l489;
  reg                 _zz_when_TxnManCS_l489_1;
  wire       [5:0]    _zz_when_TxnManCS_l489_2;
  reg        [5:0]    _zz_when_TxnManCS_l489_3;
  reg        [5:0]    _zz__zz_cntRlseReqWrRmt_0;
  wire       [7:0]    _zz_when_TxnManCS_l521;
  wire       [7:0]    _zz_when_TxnManCS_l521_1;
  wire       [11:0]   _zz_txnMem_port;
  wire       [11:0]   _zz_txnMem_port_1;
  wire       [30:0]   _zz_txnMem_port_2;
  reg                 _zz_when_TxnManCS_l621;
  wire       [31:0]   _zz_when_TxnManCS_l665;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 lkReqGetLoc_valid;
  wire                lkReqGetLoc_ready;
  wire       [0:0]    lkReqGetLoc_payload_nId;
  wire       [21:0]   lkReqGetLoc_payload_tId;
  wire       [2:0]    lkReqGetLoc_payload_tabId;
  wire       [0:0]    lkReqGetLoc_payload_snId;
  wire       [5:0]    lkReqGetLoc_payload_txnId;
  wire       [1:0]    lkReqGetLoc_payload_lkType;
  wire                lkReqGetLoc_payload_lkRelease;
  wire                lkReqGetLoc_payload_txnTimeOut;
  wire                lkReqGetLoc_payload_txnAbt;
  wire       [5:0]    lkReqGetLoc_payload_lkIdx;
  wire       [2:0]    lkReqGetLoc_payload_wLen;
  reg                 lkReqRlseLoc_valid;
  wire                lkReqRlseLoc_ready;
  wire       [0:0]    lkReqRlseLoc_payload_nId;
  wire       [21:0]   lkReqRlseLoc_payload_tId;
  wire       [2:0]    lkReqRlseLoc_payload_tabId;
  wire       [0:0]    lkReqRlseLoc_payload_snId;
  wire       [5:0]    lkReqRlseLoc_payload_txnId;
  wire       [1:0]    lkReqRlseLoc_payload_lkType;
  wire                lkReqRlseLoc_payload_lkRelease;
  wire                lkReqRlseLoc_payload_txnTimeOut;
  wire                lkReqRlseLoc_payload_txnAbt;
  wire       [5:0]    lkReqRlseLoc_payload_lkIdx;
  wire       [2:0]    lkReqRlseLoc_payload_wLen;
  reg                 lkReqGetRmt_valid;
  wire                lkReqGetRmt_ready;
  wire       [0:0]    lkReqGetRmt_payload_nId;
  wire       [21:0]   lkReqGetRmt_payload_tId;
  wire       [2:0]    lkReqGetRmt_payload_tabId;
  wire       [0:0]    lkReqGetRmt_payload_snId;
  wire       [5:0]    lkReqGetRmt_payload_txnId;
  wire       [1:0]    lkReqGetRmt_payload_lkType;
  wire                lkReqGetRmt_payload_lkRelease;
  wire                lkReqGetRmt_payload_txnTimeOut;
  wire                lkReqGetRmt_payload_txnAbt;
  wire       [5:0]    lkReqGetRmt_payload_lkIdx;
  wire       [2:0]    lkReqGetRmt_payload_wLen;
  reg                 lkReqRlseRmt_valid;
  wire                lkReqRlseRmt_ready;
  wire       [0:0]    lkReqRlseRmt_payload_nId;
  wire       [21:0]   lkReqRlseRmt_payload_tId;
  wire       [2:0]    lkReqRlseRmt_payload_tabId;
  wire       [0:0]    lkReqRlseRmt_payload_snId;
  wire       [5:0]    lkReqRlseRmt_payload_txnId;
  wire       [1:0]    lkReqRlseRmt_payload_lkType;
  wire                lkReqRlseRmt_payload_lkRelease;
  wire                lkReqRlseRmt_payload_txnTimeOut;
  wire                lkReqRlseRmt_payload_txnAbt;
  wire       [5:0]    lkReqRlseRmt_payload_lkIdx;
  wire       [2:0]    lkReqRlseRmt_payload_wLen;
  wire                streamArbiter_8_io_output_s2mPipe_valid;
  reg                 streamArbiter_8_io_output_s2mPipe_ready;
  wire       [0:0]    streamArbiter_8_io_output_s2mPipe_payload_nId;
  wire       [21:0]   streamArbiter_8_io_output_s2mPipe_payload_tId;
  wire       [2:0]    streamArbiter_8_io_output_s2mPipe_payload_tabId;
  wire       [0:0]    streamArbiter_8_io_output_s2mPipe_payload_snId;
  wire       [5:0]    streamArbiter_8_io_output_s2mPipe_payload_txnId;
  wire       [1:0]    streamArbiter_8_io_output_s2mPipe_payload_lkType;
  wire                streamArbiter_8_io_output_s2mPipe_payload_lkRelease;
  wire                streamArbiter_8_io_output_s2mPipe_payload_txnTimeOut;
  wire                streamArbiter_8_io_output_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamArbiter_8_io_output_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamArbiter_8_io_output_s2mPipe_payload_wLen;
  reg                 streamArbiter_8_io_output_rValid;
  reg        [0:0]    streamArbiter_8_io_output_rData_nId;
  reg        [21:0]   streamArbiter_8_io_output_rData_tId;
  reg        [2:0]    streamArbiter_8_io_output_rData_tabId;
  reg        [0:0]    streamArbiter_8_io_output_rData_snId;
  reg        [5:0]    streamArbiter_8_io_output_rData_txnId;
  reg        [1:0]    streamArbiter_8_io_output_rData_lkType;
  reg                 streamArbiter_8_io_output_rData_lkRelease;
  reg                 streamArbiter_8_io_output_rData_txnTimeOut;
  reg                 streamArbiter_8_io_output_rData_txnAbt;
  reg        [5:0]    streamArbiter_8_io_output_rData_lkIdx;
  reg        [2:0]    streamArbiter_8_io_output_rData_wLen;
  wire       [1:0]    _zz_payload_lkType;
  wire                streamArbiter_8_io_output_s2mPipe_m2sPipe_valid;
  wire                streamArbiter_8_io_output_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType;
  wire                streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamArbiter_8_io_output_s2mPipe_rValid;
  reg        [0:0]    streamArbiter_8_io_output_s2mPipe_rData_nId;
  reg        [21:0]   streamArbiter_8_io_output_s2mPipe_rData_tId;
  reg        [2:0]    streamArbiter_8_io_output_s2mPipe_rData_tabId;
  reg        [0:0]    streamArbiter_8_io_output_s2mPipe_rData_snId;
  reg        [5:0]    streamArbiter_8_io_output_s2mPipe_rData_txnId;
  reg        [1:0]    streamArbiter_8_io_output_s2mPipe_rData_lkType;
  reg                 streamArbiter_8_io_output_s2mPipe_rData_lkRelease;
  reg                 streamArbiter_8_io_output_s2mPipe_rData_txnTimeOut;
  reg                 streamArbiter_8_io_output_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamArbiter_8_io_output_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamArbiter_8_io_output_s2mPipe_rData_wLen;
  wire                when_Stream_l368;
  wire                streamArbiter_9_io_output_s2mPipe_valid;
  reg                 streamArbiter_9_io_output_s2mPipe_ready;
  wire       [0:0]    streamArbiter_9_io_output_s2mPipe_payload_nId;
  wire       [21:0]   streamArbiter_9_io_output_s2mPipe_payload_tId;
  wire       [2:0]    streamArbiter_9_io_output_s2mPipe_payload_tabId;
  wire       [0:0]    streamArbiter_9_io_output_s2mPipe_payload_snId;
  wire       [5:0]    streamArbiter_9_io_output_s2mPipe_payload_txnId;
  wire       [1:0]    streamArbiter_9_io_output_s2mPipe_payload_lkType;
  wire                streamArbiter_9_io_output_s2mPipe_payload_lkRelease;
  wire                streamArbiter_9_io_output_s2mPipe_payload_txnTimeOut;
  wire                streamArbiter_9_io_output_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamArbiter_9_io_output_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamArbiter_9_io_output_s2mPipe_payload_wLen;
  reg                 streamArbiter_9_io_output_rValid;
  reg        [0:0]    streamArbiter_9_io_output_rData_nId;
  reg        [21:0]   streamArbiter_9_io_output_rData_tId;
  reg        [2:0]    streamArbiter_9_io_output_rData_tabId;
  reg        [0:0]    streamArbiter_9_io_output_rData_snId;
  reg        [5:0]    streamArbiter_9_io_output_rData_txnId;
  reg        [1:0]    streamArbiter_9_io_output_rData_lkType;
  reg                 streamArbiter_9_io_output_rData_lkRelease;
  reg                 streamArbiter_9_io_output_rData_txnTimeOut;
  reg                 streamArbiter_9_io_output_rData_txnAbt;
  reg        [5:0]    streamArbiter_9_io_output_rData_lkIdx;
  reg        [2:0]    streamArbiter_9_io_output_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_1;
  wire                streamArbiter_9_io_output_s2mPipe_m2sPipe_valid;
  wire                streamArbiter_9_io_output_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType;
  wire                streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamArbiter_9_io_output_s2mPipe_rValid;
  reg        [0:0]    streamArbiter_9_io_output_s2mPipe_rData_nId;
  reg        [21:0]   streamArbiter_9_io_output_s2mPipe_rData_tId;
  reg        [2:0]    streamArbiter_9_io_output_s2mPipe_rData_tabId;
  reg        [0:0]    streamArbiter_9_io_output_s2mPipe_rData_snId;
  reg        [5:0]    streamArbiter_9_io_output_s2mPipe_rData_txnId;
  reg        [1:0]    streamArbiter_9_io_output_s2mPipe_rData_lkType;
  reg                 streamArbiter_9_io_output_s2mPipe_rData_lkRelease;
  reg                 streamArbiter_9_io_output_s2mPipe_rData_txnTimeOut;
  reg                 streamArbiter_9_io_output_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamArbiter_9_io_output_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamArbiter_9_io_output_s2mPipe_rData_wLen;
  wire                when_Stream_l368_1;
  reg        [5:0]    cntLkReqLoc_0;
  reg        [5:0]    cntLkReqLoc_1;
  reg        [5:0]    cntLkReqLoc_2;
  reg        [5:0]    cntLkReqLoc_3;
  reg        [5:0]    cntLkReqLoc_4;
  reg        [5:0]    cntLkReqLoc_5;
  reg        [5:0]    cntLkReqLoc_6;
  reg        [5:0]    cntLkReqLoc_7;
  reg        [5:0]    cntLkReqLoc_8;
  reg        [5:0]    cntLkReqLoc_9;
  reg        [5:0]    cntLkReqLoc_10;
  reg        [5:0]    cntLkReqLoc_11;
  reg        [5:0]    cntLkReqLoc_12;
  reg        [5:0]    cntLkReqLoc_13;
  reg        [5:0]    cntLkReqLoc_14;
  reg        [5:0]    cntLkReqLoc_15;
  reg        [5:0]    cntLkReqLoc_16;
  reg        [5:0]    cntLkReqLoc_17;
  reg        [5:0]    cntLkReqLoc_18;
  reg        [5:0]    cntLkReqLoc_19;
  reg        [5:0]    cntLkReqLoc_20;
  reg        [5:0]    cntLkReqLoc_21;
  reg        [5:0]    cntLkReqLoc_22;
  reg        [5:0]    cntLkReqLoc_23;
  reg        [5:0]    cntLkReqLoc_24;
  reg        [5:0]    cntLkReqLoc_25;
  reg        [5:0]    cntLkReqLoc_26;
  reg        [5:0]    cntLkReqLoc_27;
  reg        [5:0]    cntLkReqLoc_28;
  reg        [5:0]    cntLkReqLoc_29;
  reg        [5:0]    cntLkReqLoc_30;
  reg        [5:0]    cntLkReqLoc_31;
  reg        [5:0]    cntLkReqLoc_32;
  reg        [5:0]    cntLkReqLoc_33;
  reg        [5:0]    cntLkReqLoc_34;
  reg        [5:0]    cntLkReqLoc_35;
  reg        [5:0]    cntLkReqLoc_36;
  reg        [5:0]    cntLkReqLoc_37;
  reg        [5:0]    cntLkReqLoc_38;
  reg        [5:0]    cntLkReqLoc_39;
  reg        [5:0]    cntLkReqLoc_40;
  reg        [5:0]    cntLkReqLoc_41;
  reg        [5:0]    cntLkReqLoc_42;
  reg        [5:0]    cntLkReqLoc_43;
  reg        [5:0]    cntLkReqLoc_44;
  reg        [5:0]    cntLkReqLoc_45;
  reg        [5:0]    cntLkReqLoc_46;
  reg        [5:0]    cntLkReqLoc_47;
  reg        [5:0]    cntLkReqLoc_48;
  reg        [5:0]    cntLkReqLoc_49;
  reg        [5:0]    cntLkReqLoc_50;
  reg        [5:0]    cntLkReqLoc_51;
  reg        [5:0]    cntLkReqLoc_52;
  reg        [5:0]    cntLkReqLoc_53;
  reg        [5:0]    cntLkReqLoc_54;
  reg        [5:0]    cntLkReqLoc_55;
  reg        [5:0]    cntLkReqLoc_56;
  reg        [5:0]    cntLkReqLoc_57;
  reg        [5:0]    cntLkReqLoc_58;
  reg        [5:0]    cntLkReqLoc_59;
  reg        [5:0]    cntLkReqLoc_60;
  reg        [5:0]    cntLkReqLoc_61;
  reg        [5:0]    cntLkReqLoc_62;
  reg        [5:0]    cntLkReqLoc_63;
  reg        [5:0]    cntLkReqRmt_0;
  reg        [5:0]    cntLkReqRmt_1;
  reg        [5:0]    cntLkReqRmt_2;
  reg        [5:0]    cntLkReqRmt_3;
  reg        [5:0]    cntLkReqRmt_4;
  reg        [5:0]    cntLkReqRmt_5;
  reg        [5:0]    cntLkReqRmt_6;
  reg        [5:0]    cntLkReqRmt_7;
  reg        [5:0]    cntLkReqRmt_8;
  reg        [5:0]    cntLkReqRmt_9;
  reg        [5:0]    cntLkReqRmt_10;
  reg        [5:0]    cntLkReqRmt_11;
  reg        [5:0]    cntLkReqRmt_12;
  reg        [5:0]    cntLkReqRmt_13;
  reg        [5:0]    cntLkReqRmt_14;
  reg        [5:0]    cntLkReqRmt_15;
  reg        [5:0]    cntLkReqRmt_16;
  reg        [5:0]    cntLkReqRmt_17;
  reg        [5:0]    cntLkReqRmt_18;
  reg        [5:0]    cntLkReqRmt_19;
  reg        [5:0]    cntLkReqRmt_20;
  reg        [5:0]    cntLkReqRmt_21;
  reg        [5:0]    cntLkReqRmt_22;
  reg        [5:0]    cntLkReqRmt_23;
  reg        [5:0]    cntLkReqRmt_24;
  reg        [5:0]    cntLkReqRmt_25;
  reg        [5:0]    cntLkReqRmt_26;
  reg        [5:0]    cntLkReqRmt_27;
  reg        [5:0]    cntLkReqRmt_28;
  reg        [5:0]    cntLkReqRmt_29;
  reg        [5:0]    cntLkReqRmt_30;
  reg        [5:0]    cntLkReqRmt_31;
  reg        [5:0]    cntLkReqRmt_32;
  reg        [5:0]    cntLkReqRmt_33;
  reg        [5:0]    cntLkReqRmt_34;
  reg        [5:0]    cntLkReqRmt_35;
  reg        [5:0]    cntLkReqRmt_36;
  reg        [5:0]    cntLkReqRmt_37;
  reg        [5:0]    cntLkReqRmt_38;
  reg        [5:0]    cntLkReqRmt_39;
  reg        [5:0]    cntLkReqRmt_40;
  reg        [5:0]    cntLkReqRmt_41;
  reg        [5:0]    cntLkReqRmt_42;
  reg        [5:0]    cntLkReqRmt_43;
  reg        [5:0]    cntLkReqRmt_44;
  reg        [5:0]    cntLkReqRmt_45;
  reg        [5:0]    cntLkReqRmt_46;
  reg        [5:0]    cntLkReqRmt_47;
  reg        [5:0]    cntLkReqRmt_48;
  reg        [5:0]    cntLkReqRmt_49;
  reg        [5:0]    cntLkReqRmt_50;
  reg        [5:0]    cntLkReqRmt_51;
  reg        [5:0]    cntLkReqRmt_52;
  reg        [5:0]    cntLkReqRmt_53;
  reg        [5:0]    cntLkReqRmt_54;
  reg        [5:0]    cntLkReqRmt_55;
  reg        [5:0]    cntLkReqRmt_56;
  reg        [5:0]    cntLkReqRmt_57;
  reg        [5:0]    cntLkReqRmt_58;
  reg        [5:0]    cntLkReqRmt_59;
  reg        [5:0]    cntLkReqRmt_60;
  reg        [5:0]    cntLkReqRmt_61;
  reg        [5:0]    cntLkReqRmt_62;
  reg        [5:0]    cntLkReqRmt_63;
  reg        [5:0]    cntLkRespLoc_0;
  reg        [5:0]    cntLkRespLoc_1;
  reg        [5:0]    cntLkRespLoc_2;
  reg        [5:0]    cntLkRespLoc_3;
  reg        [5:0]    cntLkRespLoc_4;
  reg        [5:0]    cntLkRespLoc_5;
  reg        [5:0]    cntLkRespLoc_6;
  reg        [5:0]    cntLkRespLoc_7;
  reg        [5:0]    cntLkRespLoc_8;
  reg        [5:0]    cntLkRespLoc_9;
  reg        [5:0]    cntLkRespLoc_10;
  reg        [5:0]    cntLkRespLoc_11;
  reg        [5:0]    cntLkRespLoc_12;
  reg        [5:0]    cntLkRespLoc_13;
  reg        [5:0]    cntLkRespLoc_14;
  reg        [5:0]    cntLkRespLoc_15;
  reg        [5:0]    cntLkRespLoc_16;
  reg        [5:0]    cntLkRespLoc_17;
  reg        [5:0]    cntLkRespLoc_18;
  reg        [5:0]    cntLkRespLoc_19;
  reg        [5:0]    cntLkRespLoc_20;
  reg        [5:0]    cntLkRespLoc_21;
  reg        [5:0]    cntLkRespLoc_22;
  reg        [5:0]    cntLkRespLoc_23;
  reg        [5:0]    cntLkRespLoc_24;
  reg        [5:0]    cntLkRespLoc_25;
  reg        [5:0]    cntLkRespLoc_26;
  reg        [5:0]    cntLkRespLoc_27;
  reg        [5:0]    cntLkRespLoc_28;
  reg        [5:0]    cntLkRespLoc_29;
  reg        [5:0]    cntLkRespLoc_30;
  reg        [5:0]    cntLkRespLoc_31;
  reg        [5:0]    cntLkRespLoc_32;
  reg        [5:0]    cntLkRespLoc_33;
  reg        [5:0]    cntLkRespLoc_34;
  reg        [5:0]    cntLkRespLoc_35;
  reg        [5:0]    cntLkRespLoc_36;
  reg        [5:0]    cntLkRespLoc_37;
  reg        [5:0]    cntLkRespLoc_38;
  reg        [5:0]    cntLkRespLoc_39;
  reg        [5:0]    cntLkRespLoc_40;
  reg        [5:0]    cntLkRespLoc_41;
  reg        [5:0]    cntLkRespLoc_42;
  reg        [5:0]    cntLkRespLoc_43;
  reg        [5:0]    cntLkRespLoc_44;
  reg        [5:0]    cntLkRespLoc_45;
  reg        [5:0]    cntLkRespLoc_46;
  reg        [5:0]    cntLkRespLoc_47;
  reg        [5:0]    cntLkRespLoc_48;
  reg        [5:0]    cntLkRespLoc_49;
  reg        [5:0]    cntLkRespLoc_50;
  reg        [5:0]    cntLkRespLoc_51;
  reg        [5:0]    cntLkRespLoc_52;
  reg        [5:0]    cntLkRespLoc_53;
  reg        [5:0]    cntLkRespLoc_54;
  reg        [5:0]    cntLkRespLoc_55;
  reg        [5:0]    cntLkRespLoc_56;
  reg        [5:0]    cntLkRespLoc_57;
  reg        [5:0]    cntLkRespLoc_58;
  reg        [5:0]    cntLkRespLoc_59;
  reg        [5:0]    cntLkRespLoc_60;
  reg        [5:0]    cntLkRespLoc_61;
  reg        [5:0]    cntLkRespLoc_62;
  reg        [5:0]    cntLkRespLoc_63;
  reg        [5:0]    cntLkRespRmt_0;
  reg        [5:0]    cntLkRespRmt_1;
  reg        [5:0]    cntLkRespRmt_2;
  reg        [5:0]    cntLkRespRmt_3;
  reg        [5:0]    cntLkRespRmt_4;
  reg        [5:0]    cntLkRespRmt_5;
  reg        [5:0]    cntLkRespRmt_6;
  reg        [5:0]    cntLkRespRmt_7;
  reg        [5:0]    cntLkRespRmt_8;
  reg        [5:0]    cntLkRespRmt_9;
  reg        [5:0]    cntLkRespRmt_10;
  reg        [5:0]    cntLkRespRmt_11;
  reg        [5:0]    cntLkRespRmt_12;
  reg        [5:0]    cntLkRespRmt_13;
  reg        [5:0]    cntLkRespRmt_14;
  reg        [5:0]    cntLkRespRmt_15;
  reg        [5:0]    cntLkRespRmt_16;
  reg        [5:0]    cntLkRespRmt_17;
  reg        [5:0]    cntLkRespRmt_18;
  reg        [5:0]    cntLkRespRmt_19;
  reg        [5:0]    cntLkRespRmt_20;
  reg        [5:0]    cntLkRespRmt_21;
  reg        [5:0]    cntLkRespRmt_22;
  reg        [5:0]    cntLkRespRmt_23;
  reg        [5:0]    cntLkRespRmt_24;
  reg        [5:0]    cntLkRespRmt_25;
  reg        [5:0]    cntLkRespRmt_26;
  reg        [5:0]    cntLkRespRmt_27;
  reg        [5:0]    cntLkRespRmt_28;
  reg        [5:0]    cntLkRespRmt_29;
  reg        [5:0]    cntLkRespRmt_30;
  reg        [5:0]    cntLkRespRmt_31;
  reg        [5:0]    cntLkRespRmt_32;
  reg        [5:0]    cntLkRespRmt_33;
  reg        [5:0]    cntLkRespRmt_34;
  reg        [5:0]    cntLkRespRmt_35;
  reg        [5:0]    cntLkRespRmt_36;
  reg        [5:0]    cntLkRespRmt_37;
  reg        [5:0]    cntLkRespRmt_38;
  reg        [5:0]    cntLkRespRmt_39;
  reg        [5:0]    cntLkRespRmt_40;
  reg        [5:0]    cntLkRespRmt_41;
  reg        [5:0]    cntLkRespRmt_42;
  reg        [5:0]    cntLkRespRmt_43;
  reg        [5:0]    cntLkRespRmt_44;
  reg        [5:0]    cntLkRespRmt_45;
  reg        [5:0]    cntLkRespRmt_46;
  reg        [5:0]    cntLkRespRmt_47;
  reg        [5:0]    cntLkRespRmt_48;
  reg        [5:0]    cntLkRespRmt_49;
  reg        [5:0]    cntLkRespRmt_50;
  reg        [5:0]    cntLkRespRmt_51;
  reg        [5:0]    cntLkRespRmt_52;
  reg        [5:0]    cntLkRespRmt_53;
  reg        [5:0]    cntLkRespRmt_54;
  reg        [5:0]    cntLkRespRmt_55;
  reg        [5:0]    cntLkRespRmt_56;
  reg        [5:0]    cntLkRespRmt_57;
  reg        [5:0]    cntLkRespRmt_58;
  reg        [5:0]    cntLkRespRmt_59;
  reg        [5:0]    cntLkRespRmt_60;
  reg        [5:0]    cntLkRespRmt_61;
  reg        [5:0]    cntLkRespRmt_62;
  reg        [5:0]    cntLkRespRmt_63;
  reg        [5:0]    cntLkHoldLoc_0;
  reg        [5:0]    cntLkHoldLoc_1;
  reg        [5:0]    cntLkHoldLoc_2;
  reg        [5:0]    cntLkHoldLoc_3;
  reg        [5:0]    cntLkHoldLoc_4;
  reg        [5:0]    cntLkHoldLoc_5;
  reg        [5:0]    cntLkHoldLoc_6;
  reg        [5:0]    cntLkHoldLoc_7;
  reg        [5:0]    cntLkHoldLoc_8;
  reg        [5:0]    cntLkHoldLoc_9;
  reg        [5:0]    cntLkHoldLoc_10;
  reg        [5:0]    cntLkHoldLoc_11;
  reg        [5:0]    cntLkHoldLoc_12;
  reg        [5:0]    cntLkHoldLoc_13;
  reg        [5:0]    cntLkHoldLoc_14;
  reg        [5:0]    cntLkHoldLoc_15;
  reg        [5:0]    cntLkHoldLoc_16;
  reg        [5:0]    cntLkHoldLoc_17;
  reg        [5:0]    cntLkHoldLoc_18;
  reg        [5:0]    cntLkHoldLoc_19;
  reg        [5:0]    cntLkHoldLoc_20;
  reg        [5:0]    cntLkHoldLoc_21;
  reg        [5:0]    cntLkHoldLoc_22;
  reg        [5:0]    cntLkHoldLoc_23;
  reg        [5:0]    cntLkHoldLoc_24;
  reg        [5:0]    cntLkHoldLoc_25;
  reg        [5:0]    cntLkHoldLoc_26;
  reg        [5:0]    cntLkHoldLoc_27;
  reg        [5:0]    cntLkHoldLoc_28;
  reg        [5:0]    cntLkHoldLoc_29;
  reg        [5:0]    cntLkHoldLoc_30;
  reg        [5:0]    cntLkHoldLoc_31;
  reg        [5:0]    cntLkHoldLoc_32;
  reg        [5:0]    cntLkHoldLoc_33;
  reg        [5:0]    cntLkHoldLoc_34;
  reg        [5:0]    cntLkHoldLoc_35;
  reg        [5:0]    cntLkHoldLoc_36;
  reg        [5:0]    cntLkHoldLoc_37;
  reg        [5:0]    cntLkHoldLoc_38;
  reg        [5:0]    cntLkHoldLoc_39;
  reg        [5:0]    cntLkHoldLoc_40;
  reg        [5:0]    cntLkHoldLoc_41;
  reg        [5:0]    cntLkHoldLoc_42;
  reg        [5:0]    cntLkHoldLoc_43;
  reg        [5:0]    cntLkHoldLoc_44;
  reg        [5:0]    cntLkHoldLoc_45;
  reg        [5:0]    cntLkHoldLoc_46;
  reg        [5:0]    cntLkHoldLoc_47;
  reg        [5:0]    cntLkHoldLoc_48;
  reg        [5:0]    cntLkHoldLoc_49;
  reg        [5:0]    cntLkHoldLoc_50;
  reg        [5:0]    cntLkHoldLoc_51;
  reg        [5:0]    cntLkHoldLoc_52;
  reg        [5:0]    cntLkHoldLoc_53;
  reg        [5:0]    cntLkHoldLoc_54;
  reg        [5:0]    cntLkHoldLoc_55;
  reg        [5:0]    cntLkHoldLoc_56;
  reg        [5:0]    cntLkHoldLoc_57;
  reg        [5:0]    cntLkHoldLoc_58;
  reg        [5:0]    cntLkHoldLoc_59;
  reg        [5:0]    cntLkHoldLoc_60;
  reg        [5:0]    cntLkHoldLoc_61;
  reg        [5:0]    cntLkHoldLoc_62;
  reg        [5:0]    cntLkHoldLoc_63;
  reg        [5:0]    cntLkHoldRmt_0;
  reg        [5:0]    cntLkHoldRmt_1;
  reg        [5:0]    cntLkHoldRmt_2;
  reg        [5:0]    cntLkHoldRmt_3;
  reg        [5:0]    cntLkHoldRmt_4;
  reg        [5:0]    cntLkHoldRmt_5;
  reg        [5:0]    cntLkHoldRmt_6;
  reg        [5:0]    cntLkHoldRmt_7;
  reg        [5:0]    cntLkHoldRmt_8;
  reg        [5:0]    cntLkHoldRmt_9;
  reg        [5:0]    cntLkHoldRmt_10;
  reg        [5:0]    cntLkHoldRmt_11;
  reg        [5:0]    cntLkHoldRmt_12;
  reg        [5:0]    cntLkHoldRmt_13;
  reg        [5:0]    cntLkHoldRmt_14;
  reg        [5:0]    cntLkHoldRmt_15;
  reg        [5:0]    cntLkHoldRmt_16;
  reg        [5:0]    cntLkHoldRmt_17;
  reg        [5:0]    cntLkHoldRmt_18;
  reg        [5:0]    cntLkHoldRmt_19;
  reg        [5:0]    cntLkHoldRmt_20;
  reg        [5:0]    cntLkHoldRmt_21;
  reg        [5:0]    cntLkHoldRmt_22;
  reg        [5:0]    cntLkHoldRmt_23;
  reg        [5:0]    cntLkHoldRmt_24;
  reg        [5:0]    cntLkHoldRmt_25;
  reg        [5:0]    cntLkHoldRmt_26;
  reg        [5:0]    cntLkHoldRmt_27;
  reg        [5:0]    cntLkHoldRmt_28;
  reg        [5:0]    cntLkHoldRmt_29;
  reg        [5:0]    cntLkHoldRmt_30;
  reg        [5:0]    cntLkHoldRmt_31;
  reg        [5:0]    cntLkHoldRmt_32;
  reg        [5:0]    cntLkHoldRmt_33;
  reg        [5:0]    cntLkHoldRmt_34;
  reg        [5:0]    cntLkHoldRmt_35;
  reg        [5:0]    cntLkHoldRmt_36;
  reg        [5:0]    cntLkHoldRmt_37;
  reg        [5:0]    cntLkHoldRmt_38;
  reg        [5:0]    cntLkHoldRmt_39;
  reg        [5:0]    cntLkHoldRmt_40;
  reg        [5:0]    cntLkHoldRmt_41;
  reg        [5:0]    cntLkHoldRmt_42;
  reg        [5:0]    cntLkHoldRmt_43;
  reg        [5:0]    cntLkHoldRmt_44;
  reg        [5:0]    cntLkHoldRmt_45;
  reg        [5:0]    cntLkHoldRmt_46;
  reg        [5:0]    cntLkHoldRmt_47;
  reg        [5:0]    cntLkHoldRmt_48;
  reg        [5:0]    cntLkHoldRmt_49;
  reg        [5:0]    cntLkHoldRmt_50;
  reg        [5:0]    cntLkHoldRmt_51;
  reg        [5:0]    cntLkHoldRmt_52;
  reg        [5:0]    cntLkHoldRmt_53;
  reg        [5:0]    cntLkHoldRmt_54;
  reg        [5:0]    cntLkHoldRmt_55;
  reg        [5:0]    cntLkHoldRmt_56;
  reg        [5:0]    cntLkHoldRmt_57;
  reg        [5:0]    cntLkHoldRmt_58;
  reg        [5:0]    cntLkHoldRmt_59;
  reg        [5:0]    cntLkHoldRmt_60;
  reg        [5:0]    cntLkHoldRmt_61;
  reg        [5:0]    cntLkHoldRmt_62;
  reg        [5:0]    cntLkHoldRmt_63;
  reg        [5:0]    cntLkWaitLoc_0;
  reg        [5:0]    cntLkWaitLoc_1;
  reg        [5:0]    cntLkWaitLoc_2;
  reg        [5:0]    cntLkWaitLoc_3;
  reg        [5:0]    cntLkWaitLoc_4;
  reg        [5:0]    cntLkWaitLoc_5;
  reg        [5:0]    cntLkWaitLoc_6;
  reg        [5:0]    cntLkWaitLoc_7;
  reg        [5:0]    cntLkWaitLoc_8;
  reg        [5:0]    cntLkWaitLoc_9;
  reg        [5:0]    cntLkWaitLoc_10;
  reg        [5:0]    cntLkWaitLoc_11;
  reg        [5:0]    cntLkWaitLoc_12;
  reg        [5:0]    cntLkWaitLoc_13;
  reg        [5:0]    cntLkWaitLoc_14;
  reg        [5:0]    cntLkWaitLoc_15;
  reg        [5:0]    cntLkWaitLoc_16;
  reg        [5:0]    cntLkWaitLoc_17;
  reg        [5:0]    cntLkWaitLoc_18;
  reg        [5:0]    cntLkWaitLoc_19;
  reg        [5:0]    cntLkWaitLoc_20;
  reg        [5:0]    cntLkWaitLoc_21;
  reg        [5:0]    cntLkWaitLoc_22;
  reg        [5:0]    cntLkWaitLoc_23;
  reg        [5:0]    cntLkWaitLoc_24;
  reg        [5:0]    cntLkWaitLoc_25;
  reg        [5:0]    cntLkWaitLoc_26;
  reg        [5:0]    cntLkWaitLoc_27;
  reg        [5:0]    cntLkWaitLoc_28;
  reg        [5:0]    cntLkWaitLoc_29;
  reg        [5:0]    cntLkWaitLoc_30;
  reg        [5:0]    cntLkWaitLoc_31;
  reg        [5:0]    cntLkWaitLoc_32;
  reg        [5:0]    cntLkWaitLoc_33;
  reg        [5:0]    cntLkWaitLoc_34;
  reg        [5:0]    cntLkWaitLoc_35;
  reg        [5:0]    cntLkWaitLoc_36;
  reg        [5:0]    cntLkWaitLoc_37;
  reg        [5:0]    cntLkWaitLoc_38;
  reg        [5:0]    cntLkWaitLoc_39;
  reg        [5:0]    cntLkWaitLoc_40;
  reg        [5:0]    cntLkWaitLoc_41;
  reg        [5:0]    cntLkWaitLoc_42;
  reg        [5:0]    cntLkWaitLoc_43;
  reg        [5:0]    cntLkWaitLoc_44;
  reg        [5:0]    cntLkWaitLoc_45;
  reg        [5:0]    cntLkWaitLoc_46;
  reg        [5:0]    cntLkWaitLoc_47;
  reg        [5:0]    cntLkWaitLoc_48;
  reg        [5:0]    cntLkWaitLoc_49;
  reg        [5:0]    cntLkWaitLoc_50;
  reg        [5:0]    cntLkWaitLoc_51;
  reg        [5:0]    cntLkWaitLoc_52;
  reg        [5:0]    cntLkWaitLoc_53;
  reg        [5:0]    cntLkWaitLoc_54;
  reg        [5:0]    cntLkWaitLoc_55;
  reg        [5:0]    cntLkWaitLoc_56;
  reg        [5:0]    cntLkWaitLoc_57;
  reg        [5:0]    cntLkWaitLoc_58;
  reg        [5:0]    cntLkWaitLoc_59;
  reg        [5:0]    cntLkWaitLoc_60;
  reg        [5:0]    cntLkWaitLoc_61;
  reg        [5:0]    cntLkWaitLoc_62;
  reg        [5:0]    cntLkWaitLoc_63;
  reg        [5:0]    cntLkWaitRmt_0;
  reg        [5:0]    cntLkWaitRmt_1;
  reg        [5:0]    cntLkWaitRmt_2;
  reg        [5:0]    cntLkWaitRmt_3;
  reg        [5:0]    cntLkWaitRmt_4;
  reg        [5:0]    cntLkWaitRmt_5;
  reg        [5:0]    cntLkWaitRmt_6;
  reg        [5:0]    cntLkWaitRmt_7;
  reg        [5:0]    cntLkWaitRmt_8;
  reg        [5:0]    cntLkWaitRmt_9;
  reg        [5:0]    cntLkWaitRmt_10;
  reg        [5:0]    cntLkWaitRmt_11;
  reg        [5:0]    cntLkWaitRmt_12;
  reg        [5:0]    cntLkWaitRmt_13;
  reg        [5:0]    cntLkWaitRmt_14;
  reg        [5:0]    cntLkWaitRmt_15;
  reg        [5:0]    cntLkWaitRmt_16;
  reg        [5:0]    cntLkWaitRmt_17;
  reg        [5:0]    cntLkWaitRmt_18;
  reg        [5:0]    cntLkWaitRmt_19;
  reg        [5:0]    cntLkWaitRmt_20;
  reg        [5:0]    cntLkWaitRmt_21;
  reg        [5:0]    cntLkWaitRmt_22;
  reg        [5:0]    cntLkWaitRmt_23;
  reg        [5:0]    cntLkWaitRmt_24;
  reg        [5:0]    cntLkWaitRmt_25;
  reg        [5:0]    cntLkWaitRmt_26;
  reg        [5:0]    cntLkWaitRmt_27;
  reg        [5:0]    cntLkWaitRmt_28;
  reg        [5:0]    cntLkWaitRmt_29;
  reg        [5:0]    cntLkWaitRmt_30;
  reg        [5:0]    cntLkWaitRmt_31;
  reg        [5:0]    cntLkWaitRmt_32;
  reg        [5:0]    cntLkWaitRmt_33;
  reg        [5:0]    cntLkWaitRmt_34;
  reg        [5:0]    cntLkWaitRmt_35;
  reg        [5:0]    cntLkWaitRmt_36;
  reg        [5:0]    cntLkWaitRmt_37;
  reg        [5:0]    cntLkWaitRmt_38;
  reg        [5:0]    cntLkWaitRmt_39;
  reg        [5:0]    cntLkWaitRmt_40;
  reg        [5:0]    cntLkWaitRmt_41;
  reg        [5:0]    cntLkWaitRmt_42;
  reg        [5:0]    cntLkWaitRmt_43;
  reg        [5:0]    cntLkWaitRmt_44;
  reg        [5:0]    cntLkWaitRmt_45;
  reg        [5:0]    cntLkWaitRmt_46;
  reg        [5:0]    cntLkWaitRmt_47;
  reg        [5:0]    cntLkWaitRmt_48;
  reg        [5:0]    cntLkWaitRmt_49;
  reg        [5:0]    cntLkWaitRmt_50;
  reg        [5:0]    cntLkWaitRmt_51;
  reg        [5:0]    cntLkWaitRmt_52;
  reg        [5:0]    cntLkWaitRmt_53;
  reg        [5:0]    cntLkWaitRmt_54;
  reg        [5:0]    cntLkWaitRmt_55;
  reg        [5:0]    cntLkWaitRmt_56;
  reg        [5:0]    cntLkWaitRmt_57;
  reg        [5:0]    cntLkWaitRmt_58;
  reg        [5:0]    cntLkWaitRmt_59;
  reg        [5:0]    cntLkWaitRmt_60;
  reg        [5:0]    cntLkWaitRmt_61;
  reg        [5:0]    cntLkWaitRmt_62;
  reg        [5:0]    cntLkWaitRmt_63;
  reg        [5:0]    cntLkReqWrLoc_0;
  reg        [5:0]    cntLkReqWrLoc_1;
  reg        [5:0]    cntLkReqWrLoc_2;
  reg        [5:0]    cntLkReqWrLoc_3;
  reg        [5:0]    cntLkReqWrLoc_4;
  reg        [5:0]    cntLkReqWrLoc_5;
  reg        [5:0]    cntLkReqWrLoc_6;
  reg        [5:0]    cntLkReqWrLoc_7;
  reg        [5:0]    cntLkReqWrLoc_8;
  reg        [5:0]    cntLkReqWrLoc_9;
  reg        [5:0]    cntLkReqWrLoc_10;
  reg        [5:0]    cntLkReqWrLoc_11;
  reg        [5:0]    cntLkReqWrLoc_12;
  reg        [5:0]    cntLkReqWrLoc_13;
  reg        [5:0]    cntLkReqWrLoc_14;
  reg        [5:0]    cntLkReqWrLoc_15;
  reg        [5:0]    cntLkReqWrLoc_16;
  reg        [5:0]    cntLkReqWrLoc_17;
  reg        [5:0]    cntLkReqWrLoc_18;
  reg        [5:0]    cntLkReqWrLoc_19;
  reg        [5:0]    cntLkReqWrLoc_20;
  reg        [5:0]    cntLkReqWrLoc_21;
  reg        [5:0]    cntLkReqWrLoc_22;
  reg        [5:0]    cntLkReqWrLoc_23;
  reg        [5:0]    cntLkReqWrLoc_24;
  reg        [5:0]    cntLkReqWrLoc_25;
  reg        [5:0]    cntLkReqWrLoc_26;
  reg        [5:0]    cntLkReqWrLoc_27;
  reg        [5:0]    cntLkReqWrLoc_28;
  reg        [5:0]    cntLkReqWrLoc_29;
  reg        [5:0]    cntLkReqWrLoc_30;
  reg        [5:0]    cntLkReqWrLoc_31;
  reg        [5:0]    cntLkReqWrLoc_32;
  reg        [5:0]    cntLkReqWrLoc_33;
  reg        [5:0]    cntLkReqWrLoc_34;
  reg        [5:0]    cntLkReqWrLoc_35;
  reg        [5:0]    cntLkReqWrLoc_36;
  reg        [5:0]    cntLkReqWrLoc_37;
  reg        [5:0]    cntLkReqWrLoc_38;
  reg        [5:0]    cntLkReqWrLoc_39;
  reg        [5:0]    cntLkReqWrLoc_40;
  reg        [5:0]    cntLkReqWrLoc_41;
  reg        [5:0]    cntLkReqWrLoc_42;
  reg        [5:0]    cntLkReqWrLoc_43;
  reg        [5:0]    cntLkReqWrLoc_44;
  reg        [5:0]    cntLkReqWrLoc_45;
  reg        [5:0]    cntLkReqWrLoc_46;
  reg        [5:0]    cntLkReqWrLoc_47;
  reg        [5:0]    cntLkReqWrLoc_48;
  reg        [5:0]    cntLkReqWrLoc_49;
  reg        [5:0]    cntLkReqWrLoc_50;
  reg        [5:0]    cntLkReqWrLoc_51;
  reg        [5:0]    cntLkReqWrLoc_52;
  reg        [5:0]    cntLkReqWrLoc_53;
  reg        [5:0]    cntLkReqWrLoc_54;
  reg        [5:0]    cntLkReqWrLoc_55;
  reg        [5:0]    cntLkReqWrLoc_56;
  reg        [5:0]    cntLkReqWrLoc_57;
  reg        [5:0]    cntLkReqWrLoc_58;
  reg        [5:0]    cntLkReqWrLoc_59;
  reg        [5:0]    cntLkReqWrLoc_60;
  reg        [5:0]    cntLkReqWrLoc_61;
  reg        [5:0]    cntLkReqWrLoc_62;
  reg        [5:0]    cntLkReqWrLoc_63;
  reg        [5:0]    cntLkReqWrRmt_0;
  reg        [5:0]    cntLkReqWrRmt_1;
  reg        [5:0]    cntLkReqWrRmt_2;
  reg        [5:0]    cntLkReqWrRmt_3;
  reg        [5:0]    cntLkReqWrRmt_4;
  reg        [5:0]    cntLkReqWrRmt_5;
  reg        [5:0]    cntLkReqWrRmt_6;
  reg        [5:0]    cntLkReqWrRmt_7;
  reg        [5:0]    cntLkReqWrRmt_8;
  reg        [5:0]    cntLkReqWrRmt_9;
  reg        [5:0]    cntLkReqWrRmt_10;
  reg        [5:0]    cntLkReqWrRmt_11;
  reg        [5:0]    cntLkReqWrRmt_12;
  reg        [5:0]    cntLkReqWrRmt_13;
  reg        [5:0]    cntLkReqWrRmt_14;
  reg        [5:0]    cntLkReqWrRmt_15;
  reg        [5:0]    cntLkReqWrRmt_16;
  reg        [5:0]    cntLkReqWrRmt_17;
  reg        [5:0]    cntLkReqWrRmt_18;
  reg        [5:0]    cntLkReqWrRmt_19;
  reg        [5:0]    cntLkReqWrRmt_20;
  reg        [5:0]    cntLkReqWrRmt_21;
  reg        [5:0]    cntLkReqWrRmt_22;
  reg        [5:0]    cntLkReqWrRmt_23;
  reg        [5:0]    cntLkReqWrRmt_24;
  reg        [5:0]    cntLkReqWrRmt_25;
  reg        [5:0]    cntLkReqWrRmt_26;
  reg        [5:0]    cntLkReqWrRmt_27;
  reg        [5:0]    cntLkReqWrRmt_28;
  reg        [5:0]    cntLkReqWrRmt_29;
  reg        [5:0]    cntLkReqWrRmt_30;
  reg        [5:0]    cntLkReqWrRmt_31;
  reg        [5:0]    cntLkReqWrRmt_32;
  reg        [5:0]    cntLkReqWrRmt_33;
  reg        [5:0]    cntLkReqWrRmt_34;
  reg        [5:0]    cntLkReqWrRmt_35;
  reg        [5:0]    cntLkReqWrRmt_36;
  reg        [5:0]    cntLkReqWrRmt_37;
  reg        [5:0]    cntLkReqWrRmt_38;
  reg        [5:0]    cntLkReqWrRmt_39;
  reg        [5:0]    cntLkReqWrRmt_40;
  reg        [5:0]    cntLkReqWrRmt_41;
  reg        [5:0]    cntLkReqWrRmt_42;
  reg        [5:0]    cntLkReqWrRmt_43;
  reg        [5:0]    cntLkReqWrRmt_44;
  reg        [5:0]    cntLkReqWrRmt_45;
  reg        [5:0]    cntLkReqWrRmt_46;
  reg        [5:0]    cntLkReqWrRmt_47;
  reg        [5:0]    cntLkReqWrRmt_48;
  reg        [5:0]    cntLkReqWrRmt_49;
  reg        [5:0]    cntLkReqWrRmt_50;
  reg        [5:0]    cntLkReqWrRmt_51;
  reg        [5:0]    cntLkReqWrRmt_52;
  reg        [5:0]    cntLkReqWrRmt_53;
  reg        [5:0]    cntLkReqWrRmt_54;
  reg        [5:0]    cntLkReqWrRmt_55;
  reg        [5:0]    cntLkReqWrRmt_56;
  reg        [5:0]    cntLkReqWrRmt_57;
  reg        [5:0]    cntLkReqWrRmt_58;
  reg        [5:0]    cntLkReqWrRmt_59;
  reg        [5:0]    cntLkReqWrRmt_60;
  reg        [5:0]    cntLkReqWrRmt_61;
  reg        [5:0]    cntLkReqWrRmt_62;
  reg        [5:0]    cntLkReqWrRmt_63;
  reg        [5:0]    cntLkHoldWrLoc_0;
  reg        [5:0]    cntLkHoldWrLoc_1;
  reg        [5:0]    cntLkHoldWrLoc_2;
  reg        [5:0]    cntLkHoldWrLoc_3;
  reg        [5:0]    cntLkHoldWrLoc_4;
  reg        [5:0]    cntLkHoldWrLoc_5;
  reg        [5:0]    cntLkHoldWrLoc_6;
  reg        [5:0]    cntLkHoldWrLoc_7;
  reg        [5:0]    cntLkHoldWrLoc_8;
  reg        [5:0]    cntLkHoldWrLoc_9;
  reg        [5:0]    cntLkHoldWrLoc_10;
  reg        [5:0]    cntLkHoldWrLoc_11;
  reg        [5:0]    cntLkHoldWrLoc_12;
  reg        [5:0]    cntLkHoldWrLoc_13;
  reg        [5:0]    cntLkHoldWrLoc_14;
  reg        [5:0]    cntLkHoldWrLoc_15;
  reg        [5:0]    cntLkHoldWrLoc_16;
  reg        [5:0]    cntLkHoldWrLoc_17;
  reg        [5:0]    cntLkHoldWrLoc_18;
  reg        [5:0]    cntLkHoldWrLoc_19;
  reg        [5:0]    cntLkHoldWrLoc_20;
  reg        [5:0]    cntLkHoldWrLoc_21;
  reg        [5:0]    cntLkHoldWrLoc_22;
  reg        [5:0]    cntLkHoldWrLoc_23;
  reg        [5:0]    cntLkHoldWrLoc_24;
  reg        [5:0]    cntLkHoldWrLoc_25;
  reg        [5:0]    cntLkHoldWrLoc_26;
  reg        [5:0]    cntLkHoldWrLoc_27;
  reg        [5:0]    cntLkHoldWrLoc_28;
  reg        [5:0]    cntLkHoldWrLoc_29;
  reg        [5:0]    cntLkHoldWrLoc_30;
  reg        [5:0]    cntLkHoldWrLoc_31;
  reg        [5:0]    cntLkHoldWrLoc_32;
  reg        [5:0]    cntLkHoldWrLoc_33;
  reg        [5:0]    cntLkHoldWrLoc_34;
  reg        [5:0]    cntLkHoldWrLoc_35;
  reg        [5:0]    cntLkHoldWrLoc_36;
  reg        [5:0]    cntLkHoldWrLoc_37;
  reg        [5:0]    cntLkHoldWrLoc_38;
  reg        [5:0]    cntLkHoldWrLoc_39;
  reg        [5:0]    cntLkHoldWrLoc_40;
  reg        [5:0]    cntLkHoldWrLoc_41;
  reg        [5:0]    cntLkHoldWrLoc_42;
  reg        [5:0]    cntLkHoldWrLoc_43;
  reg        [5:0]    cntLkHoldWrLoc_44;
  reg        [5:0]    cntLkHoldWrLoc_45;
  reg        [5:0]    cntLkHoldWrLoc_46;
  reg        [5:0]    cntLkHoldWrLoc_47;
  reg        [5:0]    cntLkHoldWrLoc_48;
  reg        [5:0]    cntLkHoldWrLoc_49;
  reg        [5:0]    cntLkHoldWrLoc_50;
  reg        [5:0]    cntLkHoldWrLoc_51;
  reg        [5:0]    cntLkHoldWrLoc_52;
  reg        [5:0]    cntLkHoldWrLoc_53;
  reg        [5:0]    cntLkHoldWrLoc_54;
  reg        [5:0]    cntLkHoldWrLoc_55;
  reg        [5:0]    cntLkHoldWrLoc_56;
  reg        [5:0]    cntLkHoldWrLoc_57;
  reg        [5:0]    cntLkHoldWrLoc_58;
  reg        [5:0]    cntLkHoldWrLoc_59;
  reg        [5:0]    cntLkHoldWrLoc_60;
  reg        [5:0]    cntLkHoldWrLoc_61;
  reg        [5:0]    cntLkHoldWrLoc_62;
  reg        [5:0]    cntLkHoldWrLoc_63;
  reg        [5:0]    cntLkHoldWrRmt_0;
  reg        [5:0]    cntLkHoldWrRmt_1;
  reg        [5:0]    cntLkHoldWrRmt_2;
  reg        [5:0]    cntLkHoldWrRmt_3;
  reg        [5:0]    cntLkHoldWrRmt_4;
  reg        [5:0]    cntLkHoldWrRmt_5;
  reg        [5:0]    cntLkHoldWrRmt_6;
  reg        [5:0]    cntLkHoldWrRmt_7;
  reg        [5:0]    cntLkHoldWrRmt_8;
  reg        [5:0]    cntLkHoldWrRmt_9;
  reg        [5:0]    cntLkHoldWrRmt_10;
  reg        [5:0]    cntLkHoldWrRmt_11;
  reg        [5:0]    cntLkHoldWrRmt_12;
  reg        [5:0]    cntLkHoldWrRmt_13;
  reg        [5:0]    cntLkHoldWrRmt_14;
  reg        [5:0]    cntLkHoldWrRmt_15;
  reg        [5:0]    cntLkHoldWrRmt_16;
  reg        [5:0]    cntLkHoldWrRmt_17;
  reg        [5:0]    cntLkHoldWrRmt_18;
  reg        [5:0]    cntLkHoldWrRmt_19;
  reg        [5:0]    cntLkHoldWrRmt_20;
  reg        [5:0]    cntLkHoldWrRmt_21;
  reg        [5:0]    cntLkHoldWrRmt_22;
  reg        [5:0]    cntLkHoldWrRmt_23;
  reg        [5:0]    cntLkHoldWrRmt_24;
  reg        [5:0]    cntLkHoldWrRmt_25;
  reg        [5:0]    cntLkHoldWrRmt_26;
  reg        [5:0]    cntLkHoldWrRmt_27;
  reg        [5:0]    cntLkHoldWrRmt_28;
  reg        [5:0]    cntLkHoldWrRmt_29;
  reg        [5:0]    cntLkHoldWrRmt_30;
  reg        [5:0]    cntLkHoldWrRmt_31;
  reg        [5:0]    cntLkHoldWrRmt_32;
  reg        [5:0]    cntLkHoldWrRmt_33;
  reg        [5:0]    cntLkHoldWrRmt_34;
  reg        [5:0]    cntLkHoldWrRmt_35;
  reg        [5:0]    cntLkHoldWrRmt_36;
  reg        [5:0]    cntLkHoldWrRmt_37;
  reg        [5:0]    cntLkHoldWrRmt_38;
  reg        [5:0]    cntLkHoldWrRmt_39;
  reg        [5:0]    cntLkHoldWrRmt_40;
  reg        [5:0]    cntLkHoldWrRmt_41;
  reg        [5:0]    cntLkHoldWrRmt_42;
  reg        [5:0]    cntLkHoldWrRmt_43;
  reg        [5:0]    cntLkHoldWrRmt_44;
  reg        [5:0]    cntLkHoldWrRmt_45;
  reg        [5:0]    cntLkHoldWrRmt_46;
  reg        [5:0]    cntLkHoldWrRmt_47;
  reg        [5:0]    cntLkHoldWrRmt_48;
  reg        [5:0]    cntLkHoldWrRmt_49;
  reg        [5:0]    cntLkHoldWrRmt_50;
  reg        [5:0]    cntLkHoldWrRmt_51;
  reg        [5:0]    cntLkHoldWrRmt_52;
  reg        [5:0]    cntLkHoldWrRmt_53;
  reg        [5:0]    cntLkHoldWrRmt_54;
  reg        [5:0]    cntLkHoldWrRmt_55;
  reg        [5:0]    cntLkHoldWrRmt_56;
  reg        [5:0]    cntLkHoldWrRmt_57;
  reg        [5:0]    cntLkHoldWrRmt_58;
  reg        [5:0]    cntLkHoldWrRmt_59;
  reg        [5:0]    cntLkHoldWrRmt_60;
  reg        [5:0]    cntLkHoldWrRmt_61;
  reg        [5:0]    cntLkHoldWrRmt_62;
  reg        [5:0]    cntLkHoldWrRmt_63;
  reg        [5:0]    cntCmtReqLoc_0;
  reg        [5:0]    cntCmtReqLoc_1;
  reg        [5:0]    cntCmtReqLoc_2;
  reg        [5:0]    cntCmtReqLoc_3;
  reg        [5:0]    cntCmtReqLoc_4;
  reg        [5:0]    cntCmtReqLoc_5;
  reg        [5:0]    cntCmtReqLoc_6;
  reg        [5:0]    cntCmtReqLoc_7;
  reg        [5:0]    cntCmtReqLoc_8;
  reg        [5:0]    cntCmtReqLoc_9;
  reg        [5:0]    cntCmtReqLoc_10;
  reg        [5:0]    cntCmtReqLoc_11;
  reg        [5:0]    cntCmtReqLoc_12;
  reg        [5:0]    cntCmtReqLoc_13;
  reg        [5:0]    cntCmtReqLoc_14;
  reg        [5:0]    cntCmtReqLoc_15;
  reg        [5:0]    cntCmtReqLoc_16;
  reg        [5:0]    cntCmtReqLoc_17;
  reg        [5:0]    cntCmtReqLoc_18;
  reg        [5:0]    cntCmtReqLoc_19;
  reg        [5:0]    cntCmtReqLoc_20;
  reg        [5:0]    cntCmtReqLoc_21;
  reg        [5:0]    cntCmtReqLoc_22;
  reg        [5:0]    cntCmtReqLoc_23;
  reg        [5:0]    cntCmtReqLoc_24;
  reg        [5:0]    cntCmtReqLoc_25;
  reg        [5:0]    cntCmtReqLoc_26;
  reg        [5:0]    cntCmtReqLoc_27;
  reg        [5:0]    cntCmtReqLoc_28;
  reg        [5:0]    cntCmtReqLoc_29;
  reg        [5:0]    cntCmtReqLoc_30;
  reg        [5:0]    cntCmtReqLoc_31;
  reg        [5:0]    cntCmtReqLoc_32;
  reg        [5:0]    cntCmtReqLoc_33;
  reg        [5:0]    cntCmtReqLoc_34;
  reg        [5:0]    cntCmtReqLoc_35;
  reg        [5:0]    cntCmtReqLoc_36;
  reg        [5:0]    cntCmtReqLoc_37;
  reg        [5:0]    cntCmtReqLoc_38;
  reg        [5:0]    cntCmtReqLoc_39;
  reg        [5:0]    cntCmtReqLoc_40;
  reg        [5:0]    cntCmtReqLoc_41;
  reg        [5:0]    cntCmtReqLoc_42;
  reg        [5:0]    cntCmtReqLoc_43;
  reg        [5:0]    cntCmtReqLoc_44;
  reg        [5:0]    cntCmtReqLoc_45;
  reg        [5:0]    cntCmtReqLoc_46;
  reg        [5:0]    cntCmtReqLoc_47;
  reg        [5:0]    cntCmtReqLoc_48;
  reg        [5:0]    cntCmtReqLoc_49;
  reg        [5:0]    cntCmtReqLoc_50;
  reg        [5:0]    cntCmtReqLoc_51;
  reg        [5:0]    cntCmtReqLoc_52;
  reg        [5:0]    cntCmtReqLoc_53;
  reg        [5:0]    cntCmtReqLoc_54;
  reg        [5:0]    cntCmtReqLoc_55;
  reg        [5:0]    cntCmtReqLoc_56;
  reg        [5:0]    cntCmtReqLoc_57;
  reg        [5:0]    cntCmtReqLoc_58;
  reg        [5:0]    cntCmtReqLoc_59;
  reg        [5:0]    cntCmtReqLoc_60;
  reg        [5:0]    cntCmtReqLoc_61;
  reg        [5:0]    cntCmtReqLoc_62;
  reg        [5:0]    cntCmtReqLoc_63;
  reg        [5:0]    cntCmtReqRmt_0;
  reg        [5:0]    cntCmtReqRmt_1;
  reg        [5:0]    cntCmtReqRmt_2;
  reg        [5:0]    cntCmtReqRmt_3;
  reg        [5:0]    cntCmtReqRmt_4;
  reg        [5:0]    cntCmtReqRmt_5;
  reg        [5:0]    cntCmtReqRmt_6;
  reg        [5:0]    cntCmtReqRmt_7;
  reg        [5:0]    cntCmtReqRmt_8;
  reg        [5:0]    cntCmtReqRmt_9;
  reg        [5:0]    cntCmtReqRmt_10;
  reg        [5:0]    cntCmtReqRmt_11;
  reg        [5:0]    cntCmtReqRmt_12;
  reg        [5:0]    cntCmtReqRmt_13;
  reg        [5:0]    cntCmtReqRmt_14;
  reg        [5:0]    cntCmtReqRmt_15;
  reg        [5:0]    cntCmtReqRmt_16;
  reg        [5:0]    cntCmtReqRmt_17;
  reg        [5:0]    cntCmtReqRmt_18;
  reg        [5:0]    cntCmtReqRmt_19;
  reg        [5:0]    cntCmtReqRmt_20;
  reg        [5:0]    cntCmtReqRmt_21;
  reg        [5:0]    cntCmtReqRmt_22;
  reg        [5:0]    cntCmtReqRmt_23;
  reg        [5:0]    cntCmtReqRmt_24;
  reg        [5:0]    cntCmtReqRmt_25;
  reg        [5:0]    cntCmtReqRmt_26;
  reg        [5:0]    cntCmtReqRmt_27;
  reg        [5:0]    cntCmtReqRmt_28;
  reg        [5:0]    cntCmtReqRmt_29;
  reg        [5:0]    cntCmtReqRmt_30;
  reg        [5:0]    cntCmtReqRmt_31;
  reg        [5:0]    cntCmtReqRmt_32;
  reg        [5:0]    cntCmtReqRmt_33;
  reg        [5:0]    cntCmtReqRmt_34;
  reg        [5:0]    cntCmtReqRmt_35;
  reg        [5:0]    cntCmtReqRmt_36;
  reg        [5:0]    cntCmtReqRmt_37;
  reg        [5:0]    cntCmtReqRmt_38;
  reg        [5:0]    cntCmtReqRmt_39;
  reg        [5:0]    cntCmtReqRmt_40;
  reg        [5:0]    cntCmtReqRmt_41;
  reg        [5:0]    cntCmtReqRmt_42;
  reg        [5:0]    cntCmtReqRmt_43;
  reg        [5:0]    cntCmtReqRmt_44;
  reg        [5:0]    cntCmtReqRmt_45;
  reg        [5:0]    cntCmtReqRmt_46;
  reg        [5:0]    cntCmtReqRmt_47;
  reg        [5:0]    cntCmtReqRmt_48;
  reg        [5:0]    cntCmtReqRmt_49;
  reg        [5:0]    cntCmtReqRmt_50;
  reg        [5:0]    cntCmtReqRmt_51;
  reg        [5:0]    cntCmtReqRmt_52;
  reg        [5:0]    cntCmtReqRmt_53;
  reg        [5:0]    cntCmtReqRmt_54;
  reg        [5:0]    cntCmtReqRmt_55;
  reg        [5:0]    cntCmtReqRmt_56;
  reg        [5:0]    cntCmtReqRmt_57;
  reg        [5:0]    cntCmtReqRmt_58;
  reg        [5:0]    cntCmtReqRmt_59;
  reg        [5:0]    cntCmtReqRmt_60;
  reg        [5:0]    cntCmtReqRmt_61;
  reg        [5:0]    cntCmtReqRmt_62;
  reg        [5:0]    cntCmtReqRmt_63;
  reg        [5:0]    cntCmtRespLoc_0;
  reg        [5:0]    cntCmtRespLoc_1;
  reg        [5:0]    cntCmtRespLoc_2;
  reg        [5:0]    cntCmtRespLoc_3;
  reg        [5:0]    cntCmtRespLoc_4;
  reg        [5:0]    cntCmtRespLoc_5;
  reg        [5:0]    cntCmtRespLoc_6;
  reg        [5:0]    cntCmtRespLoc_7;
  reg        [5:0]    cntCmtRespLoc_8;
  reg        [5:0]    cntCmtRespLoc_9;
  reg        [5:0]    cntCmtRespLoc_10;
  reg        [5:0]    cntCmtRespLoc_11;
  reg        [5:0]    cntCmtRespLoc_12;
  reg        [5:0]    cntCmtRespLoc_13;
  reg        [5:0]    cntCmtRespLoc_14;
  reg        [5:0]    cntCmtRespLoc_15;
  reg        [5:0]    cntCmtRespLoc_16;
  reg        [5:0]    cntCmtRespLoc_17;
  reg        [5:0]    cntCmtRespLoc_18;
  reg        [5:0]    cntCmtRespLoc_19;
  reg        [5:0]    cntCmtRespLoc_20;
  reg        [5:0]    cntCmtRespLoc_21;
  reg        [5:0]    cntCmtRespLoc_22;
  reg        [5:0]    cntCmtRespLoc_23;
  reg        [5:0]    cntCmtRespLoc_24;
  reg        [5:0]    cntCmtRespLoc_25;
  reg        [5:0]    cntCmtRespLoc_26;
  reg        [5:0]    cntCmtRespLoc_27;
  reg        [5:0]    cntCmtRespLoc_28;
  reg        [5:0]    cntCmtRespLoc_29;
  reg        [5:0]    cntCmtRespLoc_30;
  reg        [5:0]    cntCmtRespLoc_31;
  reg        [5:0]    cntCmtRespLoc_32;
  reg        [5:0]    cntCmtRespLoc_33;
  reg        [5:0]    cntCmtRespLoc_34;
  reg        [5:0]    cntCmtRespLoc_35;
  reg        [5:0]    cntCmtRespLoc_36;
  reg        [5:0]    cntCmtRespLoc_37;
  reg        [5:0]    cntCmtRespLoc_38;
  reg        [5:0]    cntCmtRespLoc_39;
  reg        [5:0]    cntCmtRespLoc_40;
  reg        [5:0]    cntCmtRespLoc_41;
  reg        [5:0]    cntCmtRespLoc_42;
  reg        [5:0]    cntCmtRespLoc_43;
  reg        [5:0]    cntCmtRespLoc_44;
  reg        [5:0]    cntCmtRespLoc_45;
  reg        [5:0]    cntCmtRespLoc_46;
  reg        [5:0]    cntCmtRespLoc_47;
  reg        [5:0]    cntCmtRespLoc_48;
  reg        [5:0]    cntCmtRespLoc_49;
  reg        [5:0]    cntCmtRespLoc_50;
  reg        [5:0]    cntCmtRespLoc_51;
  reg        [5:0]    cntCmtRespLoc_52;
  reg        [5:0]    cntCmtRespLoc_53;
  reg        [5:0]    cntCmtRespLoc_54;
  reg        [5:0]    cntCmtRespLoc_55;
  reg        [5:0]    cntCmtRespLoc_56;
  reg        [5:0]    cntCmtRespLoc_57;
  reg        [5:0]    cntCmtRespLoc_58;
  reg        [5:0]    cntCmtRespLoc_59;
  reg        [5:0]    cntCmtRespLoc_60;
  reg        [5:0]    cntCmtRespLoc_61;
  reg        [5:0]    cntCmtRespLoc_62;
  reg        [5:0]    cntCmtRespLoc_63;
  reg        [5:0]    cntCmtRespRmt_0;
  reg        [5:0]    cntCmtRespRmt_1;
  reg        [5:0]    cntCmtRespRmt_2;
  reg        [5:0]    cntCmtRespRmt_3;
  reg        [5:0]    cntCmtRespRmt_4;
  reg        [5:0]    cntCmtRespRmt_5;
  reg        [5:0]    cntCmtRespRmt_6;
  reg        [5:0]    cntCmtRespRmt_7;
  reg        [5:0]    cntCmtRespRmt_8;
  reg        [5:0]    cntCmtRespRmt_9;
  reg        [5:0]    cntCmtRespRmt_10;
  reg        [5:0]    cntCmtRespRmt_11;
  reg        [5:0]    cntCmtRespRmt_12;
  reg        [5:0]    cntCmtRespRmt_13;
  reg        [5:0]    cntCmtRespRmt_14;
  reg        [5:0]    cntCmtRespRmt_15;
  reg        [5:0]    cntCmtRespRmt_16;
  reg        [5:0]    cntCmtRespRmt_17;
  reg        [5:0]    cntCmtRespRmt_18;
  reg        [5:0]    cntCmtRespRmt_19;
  reg        [5:0]    cntCmtRespRmt_20;
  reg        [5:0]    cntCmtRespRmt_21;
  reg        [5:0]    cntCmtRespRmt_22;
  reg        [5:0]    cntCmtRespRmt_23;
  reg        [5:0]    cntCmtRespRmt_24;
  reg        [5:0]    cntCmtRespRmt_25;
  reg        [5:0]    cntCmtRespRmt_26;
  reg        [5:0]    cntCmtRespRmt_27;
  reg        [5:0]    cntCmtRespRmt_28;
  reg        [5:0]    cntCmtRespRmt_29;
  reg        [5:0]    cntCmtRespRmt_30;
  reg        [5:0]    cntCmtRespRmt_31;
  reg        [5:0]    cntCmtRespRmt_32;
  reg        [5:0]    cntCmtRespRmt_33;
  reg        [5:0]    cntCmtRespRmt_34;
  reg        [5:0]    cntCmtRespRmt_35;
  reg        [5:0]    cntCmtRespRmt_36;
  reg        [5:0]    cntCmtRespRmt_37;
  reg        [5:0]    cntCmtRespRmt_38;
  reg        [5:0]    cntCmtRespRmt_39;
  reg        [5:0]    cntCmtRespRmt_40;
  reg        [5:0]    cntCmtRespRmt_41;
  reg        [5:0]    cntCmtRespRmt_42;
  reg        [5:0]    cntCmtRespRmt_43;
  reg        [5:0]    cntCmtRespRmt_44;
  reg        [5:0]    cntCmtRespRmt_45;
  reg        [5:0]    cntCmtRespRmt_46;
  reg        [5:0]    cntCmtRespRmt_47;
  reg        [5:0]    cntCmtRespRmt_48;
  reg        [5:0]    cntCmtRespRmt_49;
  reg        [5:0]    cntCmtRespRmt_50;
  reg        [5:0]    cntCmtRespRmt_51;
  reg        [5:0]    cntCmtRespRmt_52;
  reg        [5:0]    cntCmtRespRmt_53;
  reg        [5:0]    cntCmtRespRmt_54;
  reg        [5:0]    cntCmtRespRmt_55;
  reg        [5:0]    cntCmtRespRmt_56;
  reg        [5:0]    cntCmtRespRmt_57;
  reg        [5:0]    cntCmtRespRmt_58;
  reg        [5:0]    cntCmtRespRmt_59;
  reg        [5:0]    cntCmtRespRmt_60;
  reg        [5:0]    cntCmtRespRmt_61;
  reg        [5:0]    cntCmtRespRmt_62;
  reg        [5:0]    cntCmtRespRmt_63;
  reg        [5:0]    cntRlseReqLoc_0;
  reg        [5:0]    cntRlseReqLoc_1;
  reg        [5:0]    cntRlseReqLoc_2;
  reg        [5:0]    cntRlseReqLoc_3;
  reg        [5:0]    cntRlseReqLoc_4;
  reg        [5:0]    cntRlseReqLoc_5;
  reg        [5:0]    cntRlseReqLoc_6;
  reg        [5:0]    cntRlseReqLoc_7;
  reg        [5:0]    cntRlseReqLoc_8;
  reg        [5:0]    cntRlseReqLoc_9;
  reg        [5:0]    cntRlseReqLoc_10;
  reg        [5:0]    cntRlseReqLoc_11;
  reg        [5:0]    cntRlseReqLoc_12;
  reg        [5:0]    cntRlseReqLoc_13;
  reg        [5:0]    cntRlseReqLoc_14;
  reg        [5:0]    cntRlseReqLoc_15;
  reg        [5:0]    cntRlseReqLoc_16;
  reg        [5:0]    cntRlseReqLoc_17;
  reg        [5:0]    cntRlseReqLoc_18;
  reg        [5:0]    cntRlseReqLoc_19;
  reg        [5:0]    cntRlseReqLoc_20;
  reg        [5:0]    cntRlseReqLoc_21;
  reg        [5:0]    cntRlseReqLoc_22;
  reg        [5:0]    cntRlseReqLoc_23;
  reg        [5:0]    cntRlseReqLoc_24;
  reg        [5:0]    cntRlseReqLoc_25;
  reg        [5:0]    cntRlseReqLoc_26;
  reg        [5:0]    cntRlseReqLoc_27;
  reg        [5:0]    cntRlseReqLoc_28;
  reg        [5:0]    cntRlseReqLoc_29;
  reg        [5:0]    cntRlseReqLoc_30;
  reg        [5:0]    cntRlseReqLoc_31;
  reg        [5:0]    cntRlseReqLoc_32;
  reg        [5:0]    cntRlseReqLoc_33;
  reg        [5:0]    cntRlseReqLoc_34;
  reg        [5:0]    cntRlseReqLoc_35;
  reg        [5:0]    cntRlseReqLoc_36;
  reg        [5:0]    cntRlseReqLoc_37;
  reg        [5:0]    cntRlseReqLoc_38;
  reg        [5:0]    cntRlseReqLoc_39;
  reg        [5:0]    cntRlseReqLoc_40;
  reg        [5:0]    cntRlseReqLoc_41;
  reg        [5:0]    cntRlseReqLoc_42;
  reg        [5:0]    cntRlseReqLoc_43;
  reg        [5:0]    cntRlseReqLoc_44;
  reg        [5:0]    cntRlseReqLoc_45;
  reg        [5:0]    cntRlseReqLoc_46;
  reg        [5:0]    cntRlseReqLoc_47;
  reg        [5:0]    cntRlseReqLoc_48;
  reg        [5:0]    cntRlseReqLoc_49;
  reg        [5:0]    cntRlseReqLoc_50;
  reg        [5:0]    cntRlseReqLoc_51;
  reg        [5:0]    cntRlseReqLoc_52;
  reg        [5:0]    cntRlseReqLoc_53;
  reg        [5:0]    cntRlseReqLoc_54;
  reg        [5:0]    cntRlseReqLoc_55;
  reg        [5:0]    cntRlseReqLoc_56;
  reg        [5:0]    cntRlseReqLoc_57;
  reg        [5:0]    cntRlseReqLoc_58;
  reg        [5:0]    cntRlseReqLoc_59;
  reg        [5:0]    cntRlseReqLoc_60;
  reg        [5:0]    cntRlseReqLoc_61;
  reg        [5:0]    cntRlseReqLoc_62;
  reg        [5:0]    cntRlseReqLoc_63;
  reg        [5:0]    cntRlseReqRmt_0;
  reg        [5:0]    cntRlseReqRmt_1;
  reg        [5:0]    cntRlseReqRmt_2;
  reg        [5:0]    cntRlseReqRmt_3;
  reg        [5:0]    cntRlseReqRmt_4;
  reg        [5:0]    cntRlseReqRmt_5;
  reg        [5:0]    cntRlseReqRmt_6;
  reg        [5:0]    cntRlseReqRmt_7;
  reg        [5:0]    cntRlseReqRmt_8;
  reg        [5:0]    cntRlseReqRmt_9;
  reg        [5:0]    cntRlseReqRmt_10;
  reg        [5:0]    cntRlseReqRmt_11;
  reg        [5:0]    cntRlseReqRmt_12;
  reg        [5:0]    cntRlseReqRmt_13;
  reg        [5:0]    cntRlseReqRmt_14;
  reg        [5:0]    cntRlseReqRmt_15;
  reg        [5:0]    cntRlseReqRmt_16;
  reg        [5:0]    cntRlseReqRmt_17;
  reg        [5:0]    cntRlseReqRmt_18;
  reg        [5:0]    cntRlseReqRmt_19;
  reg        [5:0]    cntRlseReqRmt_20;
  reg        [5:0]    cntRlseReqRmt_21;
  reg        [5:0]    cntRlseReqRmt_22;
  reg        [5:0]    cntRlseReqRmt_23;
  reg        [5:0]    cntRlseReqRmt_24;
  reg        [5:0]    cntRlseReqRmt_25;
  reg        [5:0]    cntRlseReqRmt_26;
  reg        [5:0]    cntRlseReqRmt_27;
  reg        [5:0]    cntRlseReqRmt_28;
  reg        [5:0]    cntRlseReqRmt_29;
  reg        [5:0]    cntRlseReqRmt_30;
  reg        [5:0]    cntRlseReqRmt_31;
  reg        [5:0]    cntRlseReqRmt_32;
  reg        [5:0]    cntRlseReqRmt_33;
  reg        [5:0]    cntRlseReqRmt_34;
  reg        [5:0]    cntRlseReqRmt_35;
  reg        [5:0]    cntRlseReqRmt_36;
  reg        [5:0]    cntRlseReqRmt_37;
  reg        [5:0]    cntRlseReqRmt_38;
  reg        [5:0]    cntRlseReqRmt_39;
  reg        [5:0]    cntRlseReqRmt_40;
  reg        [5:0]    cntRlseReqRmt_41;
  reg        [5:0]    cntRlseReqRmt_42;
  reg        [5:0]    cntRlseReqRmt_43;
  reg        [5:0]    cntRlseReqRmt_44;
  reg        [5:0]    cntRlseReqRmt_45;
  reg        [5:0]    cntRlseReqRmt_46;
  reg        [5:0]    cntRlseReqRmt_47;
  reg        [5:0]    cntRlseReqRmt_48;
  reg        [5:0]    cntRlseReqRmt_49;
  reg        [5:0]    cntRlseReqRmt_50;
  reg        [5:0]    cntRlseReqRmt_51;
  reg        [5:0]    cntRlseReqRmt_52;
  reg        [5:0]    cntRlseReqRmt_53;
  reg        [5:0]    cntRlseReqRmt_54;
  reg        [5:0]    cntRlseReqRmt_55;
  reg        [5:0]    cntRlseReqRmt_56;
  reg        [5:0]    cntRlseReqRmt_57;
  reg        [5:0]    cntRlseReqRmt_58;
  reg        [5:0]    cntRlseReqRmt_59;
  reg        [5:0]    cntRlseReqRmt_60;
  reg        [5:0]    cntRlseReqRmt_61;
  reg        [5:0]    cntRlseReqRmt_62;
  reg        [5:0]    cntRlseReqRmt_63;
  reg        [5:0]    cntRlseReqWrLoc_0;
  reg        [5:0]    cntRlseReqWrLoc_1;
  reg        [5:0]    cntRlseReqWrLoc_2;
  reg        [5:0]    cntRlseReqWrLoc_3;
  reg        [5:0]    cntRlseReqWrLoc_4;
  reg        [5:0]    cntRlseReqWrLoc_5;
  reg        [5:0]    cntRlseReqWrLoc_6;
  reg        [5:0]    cntRlseReqWrLoc_7;
  reg        [5:0]    cntRlseReqWrLoc_8;
  reg        [5:0]    cntRlseReqWrLoc_9;
  reg        [5:0]    cntRlseReqWrLoc_10;
  reg        [5:0]    cntRlseReqWrLoc_11;
  reg        [5:0]    cntRlseReqWrLoc_12;
  reg        [5:0]    cntRlseReqWrLoc_13;
  reg        [5:0]    cntRlseReqWrLoc_14;
  reg        [5:0]    cntRlseReqWrLoc_15;
  reg        [5:0]    cntRlseReqWrLoc_16;
  reg        [5:0]    cntRlseReqWrLoc_17;
  reg        [5:0]    cntRlseReqWrLoc_18;
  reg        [5:0]    cntRlseReqWrLoc_19;
  reg        [5:0]    cntRlseReqWrLoc_20;
  reg        [5:0]    cntRlseReqWrLoc_21;
  reg        [5:0]    cntRlseReqWrLoc_22;
  reg        [5:0]    cntRlseReqWrLoc_23;
  reg        [5:0]    cntRlseReqWrLoc_24;
  reg        [5:0]    cntRlseReqWrLoc_25;
  reg        [5:0]    cntRlseReqWrLoc_26;
  reg        [5:0]    cntRlseReqWrLoc_27;
  reg        [5:0]    cntRlseReqWrLoc_28;
  reg        [5:0]    cntRlseReqWrLoc_29;
  reg        [5:0]    cntRlseReqWrLoc_30;
  reg        [5:0]    cntRlseReqWrLoc_31;
  reg        [5:0]    cntRlseReqWrLoc_32;
  reg        [5:0]    cntRlseReqWrLoc_33;
  reg        [5:0]    cntRlseReqWrLoc_34;
  reg        [5:0]    cntRlseReqWrLoc_35;
  reg        [5:0]    cntRlseReqWrLoc_36;
  reg        [5:0]    cntRlseReqWrLoc_37;
  reg        [5:0]    cntRlseReqWrLoc_38;
  reg        [5:0]    cntRlseReqWrLoc_39;
  reg        [5:0]    cntRlseReqWrLoc_40;
  reg        [5:0]    cntRlseReqWrLoc_41;
  reg        [5:0]    cntRlseReqWrLoc_42;
  reg        [5:0]    cntRlseReqWrLoc_43;
  reg        [5:0]    cntRlseReqWrLoc_44;
  reg        [5:0]    cntRlseReqWrLoc_45;
  reg        [5:0]    cntRlseReqWrLoc_46;
  reg        [5:0]    cntRlseReqWrLoc_47;
  reg        [5:0]    cntRlseReqWrLoc_48;
  reg        [5:0]    cntRlseReqWrLoc_49;
  reg        [5:0]    cntRlseReqWrLoc_50;
  reg        [5:0]    cntRlseReqWrLoc_51;
  reg        [5:0]    cntRlseReqWrLoc_52;
  reg        [5:0]    cntRlseReqWrLoc_53;
  reg        [5:0]    cntRlseReqWrLoc_54;
  reg        [5:0]    cntRlseReqWrLoc_55;
  reg        [5:0]    cntRlseReqWrLoc_56;
  reg        [5:0]    cntRlseReqWrLoc_57;
  reg        [5:0]    cntRlseReqWrLoc_58;
  reg        [5:0]    cntRlseReqWrLoc_59;
  reg        [5:0]    cntRlseReqWrLoc_60;
  reg        [5:0]    cntRlseReqWrLoc_61;
  reg        [5:0]    cntRlseReqWrLoc_62;
  reg        [5:0]    cntRlseReqWrLoc_63;
  reg        [5:0]    cntRlseReqWrRmt_0;
  reg        [5:0]    cntRlseReqWrRmt_1;
  reg        [5:0]    cntRlseReqWrRmt_2;
  reg        [5:0]    cntRlseReqWrRmt_3;
  reg        [5:0]    cntRlseReqWrRmt_4;
  reg        [5:0]    cntRlseReqWrRmt_5;
  reg        [5:0]    cntRlseReqWrRmt_6;
  reg        [5:0]    cntRlseReqWrRmt_7;
  reg        [5:0]    cntRlseReqWrRmt_8;
  reg        [5:0]    cntRlseReqWrRmt_9;
  reg        [5:0]    cntRlseReqWrRmt_10;
  reg        [5:0]    cntRlseReqWrRmt_11;
  reg        [5:0]    cntRlseReqWrRmt_12;
  reg        [5:0]    cntRlseReqWrRmt_13;
  reg        [5:0]    cntRlseReqWrRmt_14;
  reg        [5:0]    cntRlseReqWrRmt_15;
  reg        [5:0]    cntRlseReqWrRmt_16;
  reg        [5:0]    cntRlseReqWrRmt_17;
  reg        [5:0]    cntRlseReqWrRmt_18;
  reg        [5:0]    cntRlseReqWrRmt_19;
  reg        [5:0]    cntRlseReqWrRmt_20;
  reg        [5:0]    cntRlseReqWrRmt_21;
  reg        [5:0]    cntRlseReqWrRmt_22;
  reg        [5:0]    cntRlseReqWrRmt_23;
  reg        [5:0]    cntRlseReqWrRmt_24;
  reg        [5:0]    cntRlseReqWrRmt_25;
  reg        [5:0]    cntRlseReqWrRmt_26;
  reg        [5:0]    cntRlseReqWrRmt_27;
  reg        [5:0]    cntRlseReqWrRmt_28;
  reg        [5:0]    cntRlseReqWrRmt_29;
  reg        [5:0]    cntRlseReqWrRmt_30;
  reg        [5:0]    cntRlseReqWrRmt_31;
  reg        [5:0]    cntRlseReqWrRmt_32;
  reg        [5:0]    cntRlseReqWrRmt_33;
  reg        [5:0]    cntRlseReqWrRmt_34;
  reg        [5:0]    cntRlseReqWrRmt_35;
  reg        [5:0]    cntRlseReqWrRmt_36;
  reg        [5:0]    cntRlseReqWrRmt_37;
  reg        [5:0]    cntRlseReqWrRmt_38;
  reg        [5:0]    cntRlseReqWrRmt_39;
  reg        [5:0]    cntRlseReqWrRmt_40;
  reg        [5:0]    cntRlseReqWrRmt_41;
  reg        [5:0]    cntRlseReqWrRmt_42;
  reg        [5:0]    cntRlseReqWrRmt_43;
  reg        [5:0]    cntRlseReqWrRmt_44;
  reg        [5:0]    cntRlseReqWrRmt_45;
  reg        [5:0]    cntRlseReqWrRmt_46;
  reg        [5:0]    cntRlseReqWrRmt_47;
  reg        [5:0]    cntRlseReqWrRmt_48;
  reg        [5:0]    cntRlseReqWrRmt_49;
  reg        [5:0]    cntRlseReqWrRmt_50;
  reg        [5:0]    cntRlseReqWrRmt_51;
  reg        [5:0]    cntRlseReqWrRmt_52;
  reg        [5:0]    cntRlseReqWrRmt_53;
  reg        [5:0]    cntRlseReqWrRmt_54;
  reg        [5:0]    cntRlseReqWrRmt_55;
  reg        [5:0]    cntRlseReqWrRmt_56;
  reg        [5:0]    cntRlseReqWrRmt_57;
  reg        [5:0]    cntRlseReqWrRmt_58;
  reg        [5:0]    cntRlseReqWrRmt_59;
  reg        [5:0]    cntRlseReqWrRmt_60;
  reg        [5:0]    cntRlseReqWrRmt_61;
  reg        [5:0]    cntRlseReqWrRmt_62;
  reg        [5:0]    cntRlseReqWrRmt_63;
  reg        [5:0]    cntRlseRespLoc_0;
  reg        [5:0]    cntRlseRespLoc_1;
  reg        [5:0]    cntRlseRespLoc_2;
  reg        [5:0]    cntRlseRespLoc_3;
  reg        [5:0]    cntRlseRespLoc_4;
  reg        [5:0]    cntRlseRespLoc_5;
  reg        [5:0]    cntRlseRespLoc_6;
  reg        [5:0]    cntRlseRespLoc_7;
  reg        [5:0]    cntRlseRespLoc_8;
  reg        [5:0]    cntRlseRespLoc_9;
  reg        [5:0]    cntRlseRespLoc_10;
  reg        [5:0]    cntRlseRespLoc_11;
  reg        [5:0]    cntRlseRespLoc_12;
  reg        [5:0]    cntRlseRespLoc_13;
  reg        [5:0]    cntRlseRespLoc_14;
  reg        [5:0]    cntRlseRespLoc_15;
  reg        [5:0]    cntRlseRespLoc_16;
  reg        [5:0]    cntRlseRespLoc_17;
  reg        [5:0]    cntRlseRespLoc_18;
  reg        [5:0]    cntRlseRespLoc_19;
  reg        [5:0]    cntRlseRespLoc_20;
  reg        [5:0]    cntRlseRespLoc_21;
  reg        [5:0]    cntRlseRespLoc_22;
  reg        [5:0]    cntRlseRespLoc_23;
  reg        [5:0]    cntRlseRespLoc_24;
  reg        [5:0]    cntRlseRespLoc_25;
  reg        [5:0]    cntRlseRespLoc_26;
  reg        [5:0]    cntRlseRespLoc_27;
  reg        [5:0]    cntRlseRespLoc_28;
  reg        [5:0]    cntRlseRespLoc_29;
  reg        [5:0]    cntRlseRespLoc_30;
  reg        [5:0]    cntRlseRespLoc_31;
  reg        [5:0]    cntRlseRespLoc_32;
  reg        [5:0]    cntRlseRespLoc_33;
  reg        [5:0]    cntRlseRespLoc_34;
  reg        [5:0]    cntRlseRespLoc_35;
  reg        [5:0]    cntRlseRespLoc_36;
  reg        [5:0]    cntRlseRespLoc_37;
  reg        [5:0]    cntRlseRespLoc_38;
  reg        [5:0]    cntRlseRespLoc_39;
  reg        [5:0]    cntRlseRespLoc_40;
  reg        [5:0]    cntRlseRespLoc_41;
  reg        [5:0]    cntRlseRespLoc_42;
  reg        [5:0]    cntRlseRespLoc_43;
  reg        [5:0]    cntRlseRespLoc_44;
  reg        [5:0]    cntRlseRespLoc_45;
  reg        [5:0]    cntRlseRespLoc_46;
  reg        [5:0]    cntRlseRespLoc_47;
  reg        [5:0]    cntRlseRespLoc_48;
  reg        [5:0]    cntRlseRespLoc_49;
  reg        [5:0]    cntRlseRespLoc_50;
  reg        [5:0]    cntRlseRespLoc_51;
  reg        [5:0]    cntRlseRespLoc_52;
  reg        [5:0]    cntRlseRespLoc_53;
  reg        [5:0]    cntRlseRespLoc_54;
  reg        [5:0]    cntRlseRespLoc_55;
  reg        [5:0]    cntRlseRespLoc_56;
  reg        [5:0]    cntRlseRespLoc_57;
  reg        [5:0]    cntRlseRespLoc_58;
  reg        [5:0]    cntRlseRespLoc_59;
  reg        [5:0]    cntRlseRespLoc_60;
  reg        [5:0]    cntRlseRespLoc_61;
  reg        [5:0]    cntRlseRespLoc_62;
  reg        [5:0]    cntRlseRespLoc_63;
  reg        [5:0]    cntRlseRespRmt_0;
  reg        [5:0]    cntRlseRespRmt_1;
  reg        [5:0]    cntRlseRespRmt_2;
  reg        [5:0]    cntRlseRespRmt_3;
  reg        [5:0]    cntRlseRespRmt_4;
  reg        [5:0]    cntRlseRespRmt_5;
  reg        [5:0]    cntRlseRespRmt_6;
  reg        [5:0]    cntRlseRespRmt_7;
  reg        [5:0]    cntRlseRespRmt_8;
  reg        [5:0]    cntRlseRespRmt_9;
  reg        [5:0]    cntRlseRespRmt_10;
  reg        [5:0]    cntRlseRespRmt_11;
  reg        [5:0]    cntRlseRespRmt_12;
  reg        [5:0]    cntRlseRespRmt_13;
  reg        [5:0]    cntRlseRespRmt_14;
  reg        [5:0]    cntRlseRespRmt_15;
  reg        [5:0]    cntRlseRespRmt_16;
  reg        [5:0]    cntRlseRespRmt_17;
  reg        [5:0]    cntRlseRespRmt_18;
  reg        [5:0]    cntRlseRespRmt_19;
  reg        [5:0]    cntRlseRespRmt_20;
  reg        [5:0]    cntRlseRespRmt_21;
  reg        [5:0]    cntRlseRespRmt_22;
  reg        [5:0]    cntRlseRespRmt_23;
  reg        [5:0]    cntRlseRespRmt_24;
  reg        [5:0]    cntRlseRespRmt_25;
  reg        [5:0]    cntRlseRespRmt_26;
  reg        [5:0]    cntRlseRespRmt_27;
  reg        [5:0]    cntRlseRespRmt_28;
  reg        [5:0]    cntRlseRespRmt_29;
  reg        [5:0]    cntRlseRespRmt_30;
  reg        [5:0]    cntRlseRespRmt_31;
  reg        [5:0]    cntRlseRespRmt_32;
  reg        [5:0]    cntRlseRespRmt_33;
  reg        [5:0]    cntRlseRespRmt_34;
  reg        [5:0]    cntRlseRespRmt_35;
  reg        [5:0]    cntRlseRespRmt_36;
  reg        [5:0]    cntRlseRespRmt_37;
  reg        [5:0]    cntRlseRespRmt_38;
  reg        [5:0]    cntRlseRespRmt_39;
  reg        [5:0]    cntRlseRespRmt_40;
  reg        [5:0]    cntRlseRespRmt_41;
  reg        [5:0]    cntRlseRespRmt_42;
  reg        [5:0]    cntRlseRespRmt_43;
  reg        [5:0]    cntRlseRespRmt_44;
  reg        [5:0]    cntRlseRespRmt_45;
  reg        [5:0]    cntRlseRespRmt_46;
  reg        [5:0]    cntRlseRespRmt_47;
  reg        [5:0]    cntRlseRespRmt_48;
  reg        [5:0]    cntRlseRespRmt_49;
  reg        [5:0]    cntRlseRespRmt_50;
  reg        [5:0]    cntRlseRespRmt_51;
  reg        [5:0]    cntRlseRespRmt_52;
  reg        [5:0]    cntRlseRespRmt_53;
  reg        [5:0]    cntRlseRespRmt_54;
  reg        [5:0]    cntRlseRespRmt_55;
  reg        [5:0]    cntRlseRespRmt_56;
  reg        [5:0]    cntRlseRespRmt_57;
  reg        [5:0]    cntRlseRespRmt_58;
  reg        [5:0]    cntRlseRespRmt_59;
  reg        [5:0]    cntRlseRespRmt_60;
  reg        [5:0]    cntRlseRespRmt_61;
  reg        [5:0]    cntRlseRespRmt_62;
  reg        [5:0]    cntRlseRespRmt_63;
  reg        [23:0]   cntTimeOut_0;
  reg        [23:0]   cntTimeOut_1;
  reg        [23:0]   cntTimeOut_2;
  reg        [23:0]   cntTimeOut_3;
  reg        [23:0]   cntTimeOut_4;
  reg        [23:0]   cntTimeOut_5;
  reg        [23:0]   cntTimeOut_6;
  reg        [23:0]   cntTimeOut_7;
  reg        [23:0]   cntTimeOut_8;
  reg        [23:0]   cntTimeOut_9;
  reg        [23:0]   cntTimeOut_10;
  reg        [23:0]   cntTimeOut_11;
  reg        [23:0]   cntTimeOut_12;
  reg        [23:0]   cntTimeOut_13;
  reg        [23:0]   cntTimeOut_14;
  reg        [23:0]   cntTimeOut_15;
  reg        [23:0]   cntTimeOut_16;
  reg        [23:0]   cntTimeOut_17;
  reg        [23:0]   cntTimeOut_18;
  reg        [23:0]   cntTimeOut_19;
  reg        [23:0]   cntTimeOut_20;
  reg        [23:0]   cntTimeOut_21;
  reg        [23:0]   cntTimeOut_22;
  reg        [23:0]   cntTimeOut_23;
  reg        [23:0]   cntTimeOut_24;
  reg        [23:0]   cntTimeOut_25;
  reg        [23:0]   cntTimeOut_26;
  reg        [23:0]   cntTimeOut_27;
  reg        [23:0]   cntTimeOut_28;
  reg        [23:0]   cntTimeOut_29;
  reg        [23:0]   cntTimeOut_30;
  reg        [23:0]   cntTimeOut_31;
  reg        [23:0]   cntTimeOut_32;
  reg        [23:0]   cntTimeOut_33;
  reg        [23:0]   cntTimeOut_34;
  reg        [23:0]   cntTimeOut_35;
  reg        [23:0]   cntTimeOut_36;
  reg        [23:0]   cntTimeOut_37;
  reg        [23:0]   cntTimeOut_38;
  reg        [23:0]   cntTimeOut_39;
  reg        [23:0]   cntTimeOut_40;
  reg        [23:0]   cntTimeOut_41;
  reg        [23:0]   cntTimeOut_42;
  reg        [23:0]   cntTimeOut_43;
  reg        [23:0]   cntTimeOut_44;
  reg        [23:0]   cntTimeOut_45;
  reg        [23:0]   cntTimeOut_46;
  reg        [23:0]   cntTimeOut_47;
  reg        [23:0]   cntTimeOut_48;
  reg        [23:0]   cntTimeOut_49;
  reg        [23:0]   cntTimeOut_50;
  reg        [23:0]   cntTimeOut_51;
  reg        [23:0]   cntTimeOut_52;
  reg        [23:0]   cntTimeOut_53;
  reg        [23:0]   cntTimeOut_54;
  reg        [23:0]   cntTimeOut_55;
  reg        [23:0]   cntTimeOut_56;
  reg        [23:0]   cntTimeOut_57;
  reg        [23:0]   cntTimeOut_58;
  reg        [23:0]   cntTimeOut_59;
  reg        [23:0]   cntTimeOut_60;
  reg        [23:0]   cntTimeOut_61;
  reg        [23:0]   cntTimeOut_62;
  reg        [23:0]   cntTimeOut_63;
  reg                 rTimeOut_0;
  reg                 rTimeOut_1;
  reg                 rTimeOut_2;
  reg                 rTimeOut_3;
  reg                 rTimeOut_4;
  reg                 rTimeOut_5;
  reg                 rTimeOut_6;
  reg                 rTimeOut_7;
  reg                 rTimeOut_8;
  reg                 rTimeOut_9;
  reg                 rTimeOut_10;
  reg                 rTimeOut_11;
  reg                 rTimeOut_12;
  reg                 rTimeOut_13;
  reg                 rTimeOut_14;
  reg                 rTimeOut_15;
  reg                 rTimeOut_16;
  reg                 rTimeOut_17;
  reg                 rTimeOut_18;
  reg                 rTimeOut_19;
  reg                 rTimeOut_20;
  reg                 rTimeOut_21;
  reg                 rTimeOut_22;
  reg                 rTimeOut_23;
  reg                 rTimeOut_24;
  reg                 rTimeOut_25;
  reg                 rTimeOut_26;
  reg                 rTimeOut_27;
  reg                 rTimeOut_28;
  reg                 rTimeOut_29;
  reg                 rTimeOut_30;
  reg                 rTimeOut_31;
  reg                 rTimeOut_32;
  reg                 rTimeOut_33;
  reg                 rTimeOut_34;
  reg                 rTimeOut_35;
  reg                 rTimeOut_36;
  reg                 rTimeOut_37;
  reg                 rTimeOut_38;
  reg                 rTimeOut_39;
  reg                 rTimeOut_40;
  reg                 rTimeOut_41;
  reg                 rTimeOut_42;
  reg                 rTimeOut_43;
  reg                 rTimeOut_44;
  reg                 rTimeOut_45;
  reg                 rTimeOut_46;
  reg                 rTimeOut_47;
  reg                 rTimeOut_48;
  reg                 rTimeOut_49;
  reg                 rTimeOut_50;
  reg                 rTimeOut_51;
  reg                 rTimeOut_52;
  reg                 rTimeOut_53;
  reg                 rTimeOut_54;
  reg                 rTimeOut_55;
  reg                 rTimeOut_56;
  reg                 rTimeOut_57;
  reg                 rTimeOut_58;
  reg                 rTimeOut_59;
  reg                 rTimeOut_60;
  reg                 rTimeOut_61;
  reg                 rTimeOut_62;
  reg                 rTimeOut_63;
  reg                 rAbort_0;
  reg                 rAbort_1;
  reg                 rAbort_2;
  reg                 rAbort_3;
  reg                 rAbort_4;
  reg                 rAbort_5;
  reg                 rAbort_6;
  reg                 rAbort_7;
  reg                 rAbort_8;
  reg                 rAbort_9;
  reg                 rAbort_10;
  reg                 rAbort_11;
  reg                 rAbort_12;
  reg                 rAbort_13;
  reg                 rAbort_14;
  reg                 rAbort_15;
  reg                 rAbort_16;
  reg                 rAbort_17;
  reg                 rAbort_18;
  reg                 rAbort_19;
  reg                 rAbort_20;
  reg                 rAbort_21;
  reg                 rAbort_22;
  reg                 rAbort_23;
  reg                 rAbort_24;
  reg                 rAbort_25;
  reg                 rAbort_26;
  reg                 rAbort_27;
  reg                 rAbort_28;
  reg                 rAbort_29;
  reg                 rAbort_30;
  reg                 rAbort_31;
  reg                 rAbort_32;
  reg                 rAbort_33;
  reg                 rAbort_34;
  reg                 rAbort_35;
  reg                 rAbort_36;
  reg                 rAbort_37;
  reg                 rAbort_38;
  reg                 rAbort_39;
  reg                 rAbort_40;
  reg                 rAbort_41;
  reg                 rAbort_42;
  reg                 rAbort_43;
  reg                 rAbort_44;
  reg                 rAbort_45;
  reg                 rAbort_46;
  reg                 rAbort_47;
  reg                 rAbort_48;
  reg                 rAbort_49;
  reg                 rAbort_50;
  reg                 rAbort_51;
  reg                 rAbort_52;
  reg                 rAbort_53;
  reg                 rAbort_54;
  reg                 rAbort_55;
  reg                 rAbort_56;
  reg                 rAbort_57;
  reg                 rAbort_58;
  reg                 rAbort_59;
  reg                 rAbort_60;
  reg                 rAbort_61;
  reg                 rAbort_62;
  reg                 rAbort_63;
  reg                 rReqDone_0;
  reg                 rReqDone_1;
  reg                 rReqDone_2;
  reg                 rReqDone_3;
  reg                 rReqDone_4;
  reg                 rReqDone_5;
  reg                 rReqDone_6;
  reg                 rReqDone_7;
  reg                 rReqDone_8;
  reg                 rReqDone_9;
  reg                 rReqDone_10;
  reg                 rReqDone_11;
  reg                 rReqDone_12;
  reg                 rReqDone_13;
  reg                 rReqDone_14;
  reg                 rReqDone_15;
  reg                 rReqDone_16;
  reg                 rReqDone_17;
  reg                 rReqDone_18;
  reg                 rReqDone_19;
  reg                 rReqDone_20;
  reg                 rReqDone_21;
  reg                 rReqDone_22;
  reg                 rReqDone_23;
  reg                 rReqDone_24;
  reg                 rReqDone_25;
  reg                 rReqDone_26;
  reg                 rReqDone_27;
  reg                 rReqDone_28;
  reg                 rReqDone_29;
  reg                 rReqDone_30;
  reg                 rReqDone_31;
  reg                 rReqDone_32;
  reg                 rReqDone_33;
  reg                 rReqDone_34;
  reg                 rReqDone_35;
  reg                 rReqDone_36;
  reg                 rReqDone_37;
  reg                 rReqDone_38;
  reg                 rReqDone_39;
  reg                 rReqDone_40;
  reg                 rReqDone_41;
  reg                 rReqDone_42;
  reg                 rReqDone_43;
  reg                 rReqDone_44;
  reg                 rReqDone_45;
  reg                 rReqDone_46;
  reg                 rReqDone_47;
  reg                 rReqDone_48;
  reg                 rReqDone_49;
  reg                 rReqDone_50;
  reg                 rReqDone_51;
  reg                 rReqDone_52;
  reg                 rReqDone_53;
  reg                 rReqDone_54;
  reg                 rReqDone_55;
  reg                 rReqDone_56;
  reg                 rReqDone_57;
  reg                 rReqDone_58;
  reg                 rReqDone_59;
  reg                 rReqDone_60;
  reg                 rReqDone_61;
  reg                 rReqDone_62;
  reg                 rReqDone_63;
  reg                 rRlseDone_0;
  reg                 rRlseDone_1;
  reg                 rRlseDone_2;
  reg                 rRlseDone_3;
  reg                 rRlseDone_4;
  reg                 rRlseDone_5;
  reg                 rRlseDone_6;
  reg                 rRlseDone_7;
  reg                 rRlseDone_8;
  reg                 rRlseDone_9;
  reg                 rRlseDone_10;
  reg                 rRlseDone_11;
  reg                 rRlseDone_12;
  reg                 rRlseDone_13;
  reg                 rRlseDone_14;
  reg                 rRlseDone_15;
  reg                 rRlseDone_16;
  reg                 rRlseDone_17;
  reg                 rRlseDone_18;
  reg                 rRlseDone_19;
  reg                 rRlseDone_20;
  reg                 rRlseDone_21;
  reg                 rRlseDone_22;
  reg                 rRlseDone_23;
  reg                 rRlseDone_24;
  reg                 rRlseDone_25;
  reg                 rRlseDone_26;
  reg                 rRlseDone_27;
  reg                 rRlseDone_28;
  reg                 rRlseDone_29;
  reg                 rRlseDone_30;
  reg                 rRlseDone_31;
  reg                 rRlseDone_32;
  reg                 rRlseDone_33;
  reg                 rRlseDone_34;
  reg                 rRlseDone_35;
  reg                 rRlseDone_36;
  reg                 rRlseDone_37;
  reg                 rRlseDone_38;
  reg                 rRlseDone_39;
  reg                 rRlseDone_40;
  reg                 rRlseDone_41;
  reg                 rRlseDone_42;
  reg                 rRlseDone_43;
  reg                 rRlseDone_44;
  reg                 rRlseDone_45;
  reg                 rRlseDone_46;
  reg                 rRlseDone_47;
  reg                 rRlseDone_48;
  reg                 rRlseDone_49;
  reg                 rRlseDone_50;
  reg                 rRlseDone_51;
  reg                 rRlseDone_52;
  reg                 rRlseDone_53;
  reg                 rRlseDone_54;
  reg                 rRlseDone_55;
  reg                 rRlseDone_56;
  reg                 rRlseDone_57;
  reg                 rRlseDone_58;
  reg                 rRlseDone_59;
  reg                 rRlseDone_60;
  reg                 rRlseDone_61;
  reg                 rRlseDone_62;
  reg                 rRlseDone_63;
  wire                compLkReq_wantExit;
  reg                 compLkReq_wantStart;
  wire                compLkReq_wantKill;
  reg        [5:0]    compLkReq_curTxnId;
  reg                 compLkReq_txnMemRdCmd_valid;
  wire                compLkReq_txnMemRdCmd_ready;
  reg        [11:0]   compLkReq_txnMemRdCmd_payload;
  wire                compLkReq_txnMemRd_valid;
  reg                 compLkReq_txnMemRd_ready;
  wire       [0:0]    compLkReq_txnMemRd_payload_nId;
  wire       [21:0]   compLkReq_txnMemRd_payload_tId;
  wire       [2:0]    compLkReq_txnMemRd_payload_tabId;
  wire       [1:0]    compLkReq_txnMemRd_payload_lkType;
  wire       [2:0]    compLkReq_txnMemRd_payload_wLen;
  reg                 _zz_compLkReq_txnMemRd_valid;
  wire       [1:0]    _zz_compLkReq_txnMemRd_payload_lkType;
  wire       [30:0]   _zz_compLkReq_txnMemRd_payload_nId;
  wire       [1:0]    _zz_compLkReq_txnMemRd_payload_lkType_1;
  wire                compLkReq_txnMemRd_isFree;
  reg        [5:0]    compLkReq_txnLen;
  reg        [5:0]    compLkReq_reqIdx;
  wire       [11:0]   compLkReq_txnOffs;
  wire       [1:0]    _zz_lkReqGetLoc_payload_lkType;
  wire       [1:0]    _zz_lkReqGetRmt_payload_lkType;
  wire       [63:0]   compLkReq_mskTxn2Start;
  wire       [63:0]   compLkReq_mskTxn2Start_ohFirst_input;
  wire       [63:0]   compLkReq_mskTxn2Start_ohFirst_masked;
  wire       [63:0]   compLkReq_mskTxn2Start_ohFirst_value;
  wire                _zz_compLkReq_rIdxTxn2Start;
  wire                _zz_compLkReq_rIdxTxn2Start_1;
  wire                _zz_compLkReq_rIdxTxn2Start_2;
  wire                _zz_compLkReq_rIdxTxn2Start_3;
  wire                _zz_compLkReq_rIdxTxn2Start_4;
  wire                _zz_compLkReq_rIdxTxn2Start_5;
  wire                _zz_compLkReq_rIdxTxn2Start_6;
  wire                _zz_compLkReq_rIdxTxn2Start_7;
  wire                _zz_compLkReq_rIdxTxn2Start_8;
  wire                _zz_compLkReq_rIdxTxn2Start_9;
  wire                _zz_compLkReq_rIdxTxn2Start_10;
  wire                _zz_compLkReq_rIdxTxn2Start_11;
  wire                _zz_compLkReq_rIdxTxn2Start_12;
  wire                _zz_compLkReq_rIdxTxn2Start_13;
  wire                _zz_compLkReq_rIdxTxn2Start_14;
  wire                _zz_compLkReq_rIdxTxn2Start_15;
  wire                _zz_compLkReq_rIdxTxn2Start_16;
  wire                _zz_compLkReq_rIdxTxn2Start_17;
  wire                _zz_compLkReq_rIdxTxn2Start_18;
  wire                _zz_compLkReq_rIdxTxn2Start_19;
  wire                _zz_compLkReq_rIdxTxn2Start_20;
  wire                _zz_compLkReq_rIdxTxn2Start_21;
  wire                _zz_compLkReq_rIdxTxn2Start_22;
  wire                _zz_compLkReq_rIdxTxn2Start_23;
  wire                _zz_compLkReq_rIdxTxn2Start_24;
  wire                _zz_compLkReq_rIdxTxn2Start_25;
  wire                _zz_compLkReq_rIdxTxn2Start_26;
  wire                _zz_compLkReq_rIdxTxn2Start_27;
  wire                _zz_compLkReq_rIdxTxn2Start_28;
  wire                _zz_compLkReq_rIdxTxn2Start_29;
  wire                _zz_compLkReq_rIdxTxn2Start_30;
  wire                _zz_compLkReq_rIdxTxn2Start_31;
  wire                _zz_compLkReq_rIdxTxn2Start_32;
  wire                _zz_compLkReq_rIdxTxn2Start_33;
  wire                _zz_compLkReq_rIdxTxn2Start_34;
  wire                _zz_compLkReq_rIdxTxn2Start_35;
  wire                _zz_compLkReq_rIdxTxn2Start_36;
  wire                _zz_compLkReq_rIdxTxn2Start_37;
  wire                _zz_compLkReq_rIdxTxn2Start_38;
  wire                _zz_compLkReq_rIdxTxn2Start_39;
  wire                _zz_compLkReq_rIdxTxn2Start_40;
  wire                _zz_compLkReq_rIdxTxn2Start_41;
  wire                _zz_compLkReq_rIdxTxn2Start_42;
  wire                _zz_compLkReq_rIdxTxn2Start_43;
  wire                _zz_compLkReq_rIdxTxn2Start_44;
  wire                _zz_compLkReq_rIdxTxn2Start_45;
  wire                _zz_compLkReq_rIdxTxn2Start_46;
  wire                _zz_compLkReq_rIdxTxn2Start_47;
  wire                _zz_compLkReq_rIdxTxn2Start_48;
  wire                _zz_compLkReq_rIdxTxn2Start_49;
  wire                _zz_compLkReq_rIdxTxn2Start_50;
  wire                _zz_compLkReq_rIdxTxn2Start_51;
  wire                _zz_compLkReq_rIdxTxn2Start_52;
  wire                _zz_compLkReq_rIdxTxn2Start_53;
  wire                _zz_compLkReq_rIdxTxn2Start_54;
  wire                _zz_compLkReq_rIdxTxn2Start_55;
  wire                _zz_compLkReq_rIdxTxn2Start_56;
  wire                _zz_compLkReq_rIdxTxn2Start_57;
  wire                _zz_compLkReq_rIdxTxn2Start_58;
  wire                _zz_compLkReq_rIdxTxn2Start_59;
  wire                _zz_compLkReq_rIdxTxn2Start_60;
  wire                _zz_compLkReq_rIdxTxn2Start_61;
  wire                _zz_compLkReq_rIdxTxn2Start_62;
  reg        [5:0]    compLkReq_rIdxTxn2Start;
  wire                lkReqGetLoc_fire;
  wire                lkReqGetRmt_fire;
  wire                compLkReq_lkReqFire;
  wire                compLkReq_isLocal;
  wire                compLkRespLoc_wantExit;
  reg                 compLkRespLoc_wantStart;
  wire                compLkRespLoc_wantKill;
  wire                io_lkRespLoc_fire;
  reg                 compLkRespLoc_rLkResp_valid;
  reg                 compLkRespLoc_rLkResp_ready;
  reg        [0:0]    compLkRespLoc_rLkResp_payload_nId;
  reg        [21:0]   compLkRespLoc_rLkResp_payload_tId;
  reg        [2:0]    compLkRespLoc_rLkResp_payload_tabId;
  reg        [0:0]    compLkRespLoc_rLkResp_payload_snId;
  reg        [5:0]    compLkRespLoc_rLkResp_payload_txnId;
  reg        [1:0]    compLkRespLoc_rLkResp_payload_lkType;
  reg                 compLkRespLoc_rLkResp_payload_lkRelease;
  reg                 compLkRespLoc_rLkResp_payload_txnAbt;
  reg        [5:0]    compLkRespLoc_rLkResp_payload_lkIdx;
  reg        [2:0]    compLkRespLoc_rLkResp_payload_wLen;
  reg        [1:0]    compLkRespLoc_rLkResp_payload_respType;
  reg                 compLkRespLoc_rLkResp_payload_lkWaited;
  wire       [11:0]   compLkRespLoc_txnOffs;
  wire                io_lkRespLoc_fire_1;
  reg        [5:0]    compLkRespLoc_rCurTxnId;
  wire                compLkRespLoc_getAllRlse;
  wire                compLkRespLoc_getAllLkResp;
  wire       [5:0]    _zz_cntRlseRespLoc_0;
  wire       [63:0]   _zz_5;
  wire       [5:0]    _zz_cntLkHoldLoc_0;
  wire       [63:0]   _zz_6;
  wire       [5:0]    _zz_cntLkWaitLoc_0;
  wire       [63:0]   _zz_7;
  wire                compLkRespLoc_getAllRlseTimeOut;
  wire                when_TxnManCS_l166;
  wire                io_lkReqLoc_fire;
  wire                io_lkReqRmt_fire;
  wire                compLkRespLoc_firstReqAbt;
  wire                io_lkRespLoc_fire_2;
  reg                 compLkRespLoc_rFire;
  wire                when_TxnManCS_l164;
  wire       [63:0]   _zz_8;
  wire                compLkRespRmt_wantExit;
  reg                 compLkRespRmt_wantStart;
  wire                compLkRespRmt_wantKill;
  wire                io_lkRespRmt_fire;
  reg                 compLkRespRmt_rLkResp_valid;
  reg                 compLkRespRmt_rLkResp_ready;
  reg        [0:0]    compLkRespRmt_rLkResp_payload_nId;
  reg        [21:0]   compLkRespRmt_rLkResp_payload_tId;
  reg        [2:0]    compLkRespRmt_rLkResp_payload_tabId;
  reg        [0:0]    compLkRespRmt_rLkResp_payload_snId;
  reg        [5:0]    compLkRespRmt_rLkResp_payload_txnId;
  reg        [1:0]    compLkRespRmt_rLkResp_payload_lkType;
  reg                 compLkRespRmt_rLkResp_payload_lkRelease;
  reg                 compLkRespRmt_rLkResp_payload_txnAbt;
  reg        [5:0]    compLkRespRmt_rLkResp_payload_lkIdx;
  reg        [2:0]    compLkRespRmt_rLkResp_payload_wLen;
  reg        [1:0]    compLkRespRmt_rLkResp_payload_respType;
  reg                 compLkRespRmt_rLkResp_payload_lkWaited;
  reg        [7:0]    compLkRespRmt_nBeat;
  wire       [11:0]   compLkRespRmt_txnOffs;
  wire                io_lkRespRmt_fire_1;
  reg        [5:0]    compLkRespRmt_rCurTxnId;
  wire                compLkRespRmt_getAllRlse;
  wire                compLkRespRmt_getAllLkResp;
  wire       [5:0]    _zz_cntRlseRespRmt_0;
  wire       [63:0]   _zz_9;
  wire       [5:0]    _zz_cntLkHoldRmt_0;
  wire       [63:0]   _zz_10;
  wire       [5:0]    _zz_cntLkWaitRmt_0;
  wire       [63:0]   _zz_11;
  wire                compLkRespRmt_getAllRlseTimeOut;
  wire                when_TxnManCS_l261;
  wire                io_lkReqLoc_fire_1;
  wire                io_lkReqRmt_fire_1;
  wire                compLkRespRmt_firstReqAbt;
  wire                io_lkRespRmt_fire_2;
  reg                 compLkRespRmt_rFire;
  wire                when_TxnManCS_l259;
  wire       [63:0]   _zz_12;
  wire                io_axi_b_fire;
  reg                 compAxiResp_rAxiBFire;
  reg        [5:0]    compAxiResp_rAxiBId;
  wire       [63:0]   _zz_13;
  wire       [5:0]    _zz_cntCmtRespLoc_0;
  wire                compTxnCmtLoc_wantExit;
  reg                 compTxnCmtLoc_wantStart;
  wire                compTxnCmtLoc_wantKill;
  reg        [5:0]    compTxnCmtLoc_curTxnId;
  wire       [11:0]   compTxnCmtLoc_txnOffs;
  wire       [5:0]    _zz_cntCmtReqLoc_0;
  wire       [63:0]   _zz_14;
  wire       [11:0]   _zz_compTxnCmtLoc_cmtTxn_nId;
  wire       [0:0]    compTxnCmtLoc_cmtTxn_nId;
  wire       [21:0]   compTxnCmtLoc_cmtTxn_tId;
  wire       [2:0]    compTxnCmtLoc_cmtTxn_tabId;
  wire       [1:0]    compTxnCmtLoc_cmtTxn_lkType;
  wire       [2:0]    compTxnCmtLoc_cmtTxn_wLen;
  wire       [30:0]   _zz_compTxnCmtLoc_cmtTxn_nId_1;
  wire       [1:0]    _zz_compTxnCmtLoc_cmtTxn_lkType;
  reg        [0:0]    compTxnCmtLoc_rCmtTxn_nId;
  reg        [21:0]   compTxnCmtLoc_rCmtTxn_tId;
  reg        [2:0]    compTxnCmtLoc_rCmtTxn_tabId;
  reg        [1:0]    compTxnCmtLoc_rCmtTxn_lkType;
  reg        [2:0]    compTxnCmtLoc_rCmtTxn_wLen;
  reg        [7:0]    compTxnCmtLoc_nBeat;
  wire                compTxnCmtLoc_getAllLkResp;
  wire                compLkRlseLoc_wantExit;
  reg                 compLkRlseLoc_wantStart;
  wire                compLkRlseLoc_wantKill;
  reg        [5:0]    compLkRlseLoc_curTxnId;
  wire       [11:0]   compLkRlseLoc_txnOffs;
  wire       [5:0]    _zz_cntRlseReqLoc_0;
  wire       [63:0]   _zz_15;
  wire       [11:0]   _zz_compLkRlseLoc_lkItem_nId;
  wire       [0:0]    compLkRlseLoc_lkItem_nId;
  wire       [21:0]   compLkRlseLoc_lkItem_tId;
  wire       [2:0]    compLkRlseLoc_lkItem_tabId;
  wire       [0:0]    compLkRlseLoc_lkItem_snId;
  wire       [5:0]    compLkRlseLoc_lkItem_txnId;
  wire       [1:0]    compLkRlseLoc_lkItem_lkType;
  wire                compLkRlseLoc_lkItem_lkRelease;
  wire                compLkRlseLoc_lkItem_txnAbt;
  wire       [5:0]    compLkRlseLoc_lkItem_lkIdx;
  wire       [2:0]    compLkRlseLoc_lkItem_wLen;
  wire       [1:0]    compLkRlseLoc_lkItem_respType;
  wire                compLkRlseLoc_lkItem_lkWaited;
  wire       [48:0]   _zz_compLkRlseLoc_lkItem_nId_1;
  wire       [1:0]    _zz_compLkRlseLoc_lkItem_lkType;
  wire       [1:0]    _zz_compLkRlseLoc_lkItem_respType;
  wire                compLkRlseLoc_getAllLkResp;
  wire                _zz_lkReqRlseLoc_payload_txnAbt;
  wire                _zz_lkReqRlseLoc_payload_txnTimeOut;
  wire       [1:0]    _zz_lkReqRlseLoc_payload_lkType;
  reg                 _zz_lkReqRlseLoc_payload_lkRelease;
  wire                _zz_lkReqRlseLoc_payload_txnTimeOut_1;
  reg                 _zz_lkReqRlseLoc_payload_txnAbt_1;
  reg        [5:0]    _zz_lkReqRlseLoc_payload_lkIdx;
  wire                compLkRlseRmt_wantExit;
  reg                 compLkRlseRmt_wantStart;
  wire                compLkRlseRmt_wantKill;
  reg        [5:0]    compLkRlseRmt_curTxnId;
  reg        [7:0]    compLkRlseRmt_nBeat;
  wire       [11:0]   compLkRlseRmt_txnOffs;
  wire       [5:0]    _zz_cntRlseReqRmt_0;
  wire       [63:0]   _zz_16;
  wire                _zz_17;
  wire                _zz_18;
  wire                _zz_19;
  wire                _zz_20;
  wire                _zz_21;
  wire                _zz_22;
  wire                _zz_23;
  wire                _zz_24;
  wire                _zz_25;
  wire                _zz_26;
  wire                _zz_27;
  wire                _zz_28;
  wire                _zz_29;
  wire                _zz_30;
  wire                _zz_31;
  wire                _zz_32;
  wire                _zz_33;
  wire                _zz_34;
  wire                _zz_35;
  wire                _zz_36;
  wire                _zz_37;
  wire                _zz_38;
  wire                _zz_39;
  wire                _zz_40;
  wire                _zz_41;
  wire                _zz_42;
  wire                _zz_43;
  wire                _zz_44;
  wire                _zz_45;
  wire                _zz_46;
  wire                _zz_47;
  wire                _zz_48;
  wire                _zz_49;
  wire                _zz_50;
  wire                _zz_51;
  wire                _zz_52;
  wire                _zz_53;
  wire                _zz_54;
  wire                _zz_55;
  wire                _zz_56;
  wire                _zz_57;
  wire                _zz_58;
  wire                _zz_59;
  wire                _zz_60;
  wire                _zz_61;
  wire                _zz_62;
  wire                _zz_63;
  wire                _zz_64;
  wire                _zz_65;
  wire                _zz_66;
  wire                _zz_67;
  wire                _zz_68;
  wire                _zz_69;
  wire                _zz_70;
  wire                _zz_71;
  wire                _zz_72;
  wire                _zz_73;
  wire                _zz_74;
  wire                _zz_75;
  wire                _zz_76;
  wire                _zz_77;
  wire                _zz_78;
  wire                _zz_79;
  wire                _zz_80;
  wire       [11:0]   _zz_compLkRlseRmt_lkItem_nId;
  wire       [0:0]    compLkRlseRmt_lkItem_nId;
  wire       [21:0]   compLkRlseRmt_lkItem_tId;
  wire       [2:0]    compLkRlseRmt_lkItem_tabId;
  wire       [0:0]    compLkRlseRmt_lkItem_snId;
  wire       [5:0]    compLkRlseRmt_lkItem_txnId;
  wire       [1:0]    compLkRlseRmt_lkItem_lkType;
  wire                compLkRlseRmt_lkItem_lkRelease;
  wire                compLkRlseRmt_lkItem_txnAbt;
  wire       [5:0]    compLkRlseRmt_lkItem_lkIdx;
  wire       [2:0]    compLkRlseRmt_lkItem_wLen;
  wire       [1:0]    compLkRlseRmt_lkItem_respType;
  wire                compLkRlseRmt_lkItem_lkWaited;
  wire       [48:0]   _zz_compLkRlseRmt_lkItem_nId_1;
  wire       [1:0]    _zz_compLkRlseRmt_lkItem_lkType;
  wire       [1:0]    _zz_compLkRlseRmt_lkItem_respType;
  wire                compLkRlseRmt_getAllLkResp;
  wire                _zz_lkReqRlseRmt_payload_txnAbt;
  wire                _zz_lkReqRlseRmt_payload_txnTimeOut;
  wire       [1:0]    _zz_lkReqRlseRmt_payload_lkType;
  reg                 _zz_lkReqRlseRmt_payload_lkRelease;
  wire                _zz_lkReqRlseRmt_payload_txnTimeOut_1;
  reg                 _zz_lkReqRlseRmt_payload_txnAbt_1;
  reg        [5:0]    _zz_lkReqRlseRmt_payload_lkIdx;
  wire                compTimeOut_wantExit;
  reg                 compTimeOut_wantStart;
  wire                compTimeOut_wantKill;
  wire                compLoadTxn_wantExit;
  reg                 compLoadTxn_wantStart;
  wire                compLoadTxn_wantKill;
  reg        [5:0]    compLoadTxn_curTxnId;
  reg        [31:0]   compLoadTxn_cntTxn;
  wire       [11:0]   compLoadTxn_txnOffs;
  wire                io_cmdAxi_r_fire;
  reg        [511:0]  compLoadTxn_rCmdAxiData;
  wire                io_cmdAxi_r_fire_1;
  reg                 compLoadTxn_rCmdAxiFire;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_0;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_1;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_2;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_3;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_4;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_5;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_6;
  wire       [63:0]   compLoadTxn_cmdAxiDataSlice_7;
  reg                 compLoadTxn_rTxnMemLd;
  reg                 compLoadTxn_cntTxnWordInLine_willIncrement;
  reg                 compLoadTxn_cntTxnWordInLine_willClear;
  reg        [2:0]    compLoadTxn_cntTxnWordInLine_valueNext;
  reg        [2:0]    compLoadTxn_cntTxnWordInLine_value;
  wire                compLoadTxn_cntTxnWordInLine_willOverflowIfInc;
  wire                compLoadTxn_cntTxnWordInLine_willOverflow;
  reg                 compLoadTxn_cntTxnWord_willIncrement;
  reg                 compLoadTxn_cntTxnWord_willClear;
  reg        [5:0]    compLoadTxn_cntTxnWord_valueNext;
  reg        [5:0]    compLoadTxn_cntTxnWord_value;
  wire                compLoadTxn_cntTxnWord_willOverflowIfInc;
  wire                compLoadTxn_cntTxnWord_willOverflow;
  wire       [63:0]   compLoadTxn_bitsBuff;
  wire       [30:0]   compLoadTxn_txnBuff;
  wire                when_TxnManCS_l672;
  wire                clkCnt_wantExit;
  reg                 clkCnt_wantStart;
  wire                clkCnt_wantKill;
  reg        [1:0]    compLkReq_stateReg;
  reg        [1:0]    compLkReq_stateNext;
  reg                 _zz_81;
  wire                compLkReq_txnMemRd_fire;
  wire       [11:0]   _zz_compLkReq_txnMemRdCmd_payload;
  wire       [63:0]   _zz_82;
  wire       [5:0]    _zz_cntLkReqLoc_0;
  wire       [63:0]   _zz_83;
  wire       [5:0]    _zz_cntLkReqRmt_0;
  wire                when_TxnManCS_l106;
  wire       [5:0]    _zz_cntLkReqWrLoc_0;
  wire       [63:0]   _zz_84;
  wire       [5:0]    _zz_cntLkReqWrLoc_0_1;
  wire       [5:0]    _zz_cntLkReqWrRmt_0;
  wire       [63:0]   _zz_85;
  wire       [5:0]    _zz_cntLkReqWrRmt_0_1;
  wire                when_TxnManCS_l128;
  wire       [63:0]   _zz_86;
  reg        [1:0]    compLkRespLoc_stateReg;
  reg        [1:0]    compLkRespLoc_stateNext;
  wire                io_lkRespLoc_fire_3;
  wire       [5:0]    _zz_cntLkRespLoc_0;
  wire       [63:0]   _zz_87;
  wire                _zz_88;
  wire                _zz_89;
  wire                _zz_90;
  wire                _zz_91;
  wire                _zz_92;
  wire                _zz_93;
  wire                _zz_94;
  wire                _zz_95;
  wire                _zz_96;
  wire                _zz_97;
  wire                _zz_98;
  wire                _zz_99;
  wire                _zz_100;
  wire                _zz_101;
  wire                _zz_102;
  wire                _zz_103;
  wire                _zz_104;
  wire                _zz_105;
  wire                _zz_106;
  wire                _zz_107;
  wire                _zz_108;
  wire                _zz_109;
  wire                _zz_110;
  wire                _zz_111;
  wire                _zz_112;
  wire                _zz_113;
  wire                _zz_114;
  wire                _zz_115;
  wire                _zz_116;
  wire                _zz_117;
  wire                _zz_118;
  wire                _zz_119;
  wire                _zz_120;
  wire                _zz_121;
  wire                _zz_122;
  wire                _zz_123;
  wire                _zz_124;
  wire                _zz_125;
  wire                _zz_126;
  wire                _zz_127;
  wire                _zz_128;
  wire                _zz_129;
  wire                _zz_130;
  wire                _zz_131;
  wire                _zz_132;
  wire                _zz_133;
  wire                _zz_134;
  wire                _zz_135;
  wire                _zz_136;
  wire                _zz_137;
  wire                _zz_138;
  wire                _zz_139;
  wire                _zz_140;
  wire                _zz_141;
  wire                _zz_142;
  wire                _zz_143;
  wire                _zz_144;
  wire                _zz_145;
  wire                _zz_146;
  wire                _zz_147;
  wire                _zz_148;
  wire                _zz_149;
  wire                _zz_150;
  wire                _zz_151;
  wire       [5:0]    _zz_cntLkRespLoc_0_1;
  wire                when_TxnManCS_l179;
  wire       [5:0]    _zz_cntLkHoldLoc_0_1;
  wire       [5:0]    _zz_cntLkHoldWrLoc_0;
  wire       [63:0]   _zz_152;
  wire                _zz_153;
  wire                _zz_154;
  wire                _zz_155;
  wire                _zz_156;
  wire                _zz_157;
  wire                _zz_158;
  wire                _zz_159;
  wire                _zz_160;
  wire                _zz_161;
  wire                _zz_162;
  wire                _zz_163;
  wire                _zz_164;
  wire                _zz_165;
  wire                _zz_166;
  wire                _zz_167;
  wire                _zz_168;
  wire                _zz_169;
  wire                _zz_170;
  wire                _zz_171;
  wire                _zz_172;
  wire                _zz_173;
  wire                _zz_174;
  wire                _zz_175;
  wire                _zz_176;
  wire                _zz_177;
  wire                _zz_178;
  wire                _zz_179;
  wire                _zz_180;
  wire                _zz_181;
  wire                _zz_182;
  wire                _zz_183;
  wire                _zz_184;
  wire                _zz_185;
  wire                _zz_186;
  wire                _zz_187;
  wire                _zz_188;
  wire                _zz_189;
  wire                _zz_190;
  wire                _zz_191;
  wire                _zz_192;
  wire                _zz_193;
  wire                _zz_194;
  wire                _zz_195;
  wire                _zz_196;
  wire                _zz_197;
  wire                _zz_198;
  wire                _zz_199;
  wire                _zz_200;
  wire                _zz_201;
  wire                _zz_202;
  wire                _zz_203;
  wire                _zz_204;
  wire                _zz_205;
  wire                _zz_206;
  wire                _zz_207;
  wire                _zz_208;
  wire                _zz_209;
  wire                _zz_210;
  wire                _zz_211;
  wire                _zz_212;
  wire                _zz_213;
  wire                _zz_214;
  wire                _zz_215;
  wire                _zz_216;
  wire       [5:0]    _zz_cntLkHoldWrLoc_0_1;
  wire       [5:0]    _zz_cntLkHoldWrLoc_0_2;
  wire       [5:0]    _zz_cntLkWaitLoc_0_1;
  wire       [63:0]   _zz_217;
  wire       [5:0]    _zz_cntLkRespLoc_0_2;
  wire       [5:0]    _zz_cntRlseRespLoc_0_1;
  wire                when_TxnManCS_l214;
  wire                io_axi_ar_fire;
  reg        [1:0]    compLkRespRmt_stateReg;
  reg        [1:0]    compLkRespRmt_stateNext;
  wire                io_lkRespRmt_fire_3;
  wire       [5:0]    _zz_cntLkRespRmt_0;
  wire       [63:0]   _zz_218;
  wire                _zz_219;
  wire                _zz_220;
  wire                _zz_221;
  wire                _zz_222;
  wire                _zz_223;
  wire                _zz_224;
  wire                _zz_225;
  wire                _zz_226;
  wire                _zz_227;
  wire                _zz_228;
  wire                _zz_229;
  wire                _zz_230;
  wire                _zz_231;
  wire                _zz_232;
  wire                _zz_233;
  wire                _zz_234;
  wire                _zz_235;
  wire                _zz_236;
  wire                _zz_237;
  wire                _zz_238;
  wire                _zz_239;
  wire                _zz_240;
  wire                _zz_241;
  wire                _zz_242;
  wire                _zz_243;
  wire                _zz_244;
  wire                _zz_245;
  wire                _zz_246;
  wire                _zz_247;
  wire                _zz_248;
  wire                _zz_249;
  wire                _zz_250;
  wire                _zz_251;
  wire                _zz_252;
  wire                _zz_253;
  wire                _zz_254;
  wire                _zz_255;
  wire                _zz_256;
  wire                _zz_257;
  wire                _zz_258;
  wire                _zz_259;
  wire                _zz_260;
  wire                _zz_261;
  wire                _zz_262;
  wire                _zz_263;
  wire                _zz_264;
  wire                _zz_265;
  wire                _zz_266;
  wire                _zz_267;
  wire                _zz_268;
  wire                _zz_269;
  wire                _zz_270;
  wire                _zz_271;
  wire                _zz_272;
  wire                _zz_273;
  wire                _zz_274;
  wire                _zz_275;
  wire                _zz_276;
  wire                _zz_277;
  wire                _zz_278;
  wire                _zz_279;
  wire                _zz_280;
  wire                _zz_281;
  wire                _zz_282;
  wire       [5:0]    _zz_cntLkRespRmt_0_1;
  wire                when_TxnManCS_l272;
  wire       [5:0]    _zz_cntLkHoldRmt_0_1;
  wire       [5:0]    _zz_cntLkHoldWrRmt_0;
  wire       [63:0]   _zz_283;
  wire                _zz_284;
  wire                _zz_285;
  wire                _zz_286;
  wire                _zz_287;
  wire                _zz_288;
  wire                _zz_289;
  wire                _zz_290;
  wire                _zz_291;
  wire                _zz_292;
  wire                _zz_293;
  wire                _zz_294;
  wire                _zz_295;
  wire                _zz_296;
  wire                _zz_297;
  wire                _zz_298;
  wire                _zz_299;
  wire                _zz_300;
  wire                _zz_301;
  wire                _zz_302;
  wire                _zz_303;
  wire                _zz_304;
  wire                _zz_305;
  wire                _zz_306;
  wire                _zz_307;
  wire                _zz_308;
  wire                _zz_309;
  wire                _zz_310;
  wire                _zz_311;
  wire                _zz_312;
  wire                _zz_313;
  wire                _zz_314;
  wire                _zz_315;
  wire                _zz_316;
  wire                _zz_317;
  wire                _zz_318;
  wire                _zz_319;
  wire                _zz_320;
  wire                _zz_321;
  wire                _zz_322;
  wire                _zz_323;
  wire                _zz_324;
  wire                _zz_325;
  wire                _zz_326;
  wire                _zz_327;
  wire                _zz_328;
  wire                _zz_329;
  wire                _zz_330;
  wire                _zz_331;
  wire                _zz_332;
  wire                _zz_333;
  wire                _zz_334;
  wire                _zz_335;
  wire                _zz_336;
  wire                _zz_337;
  wire                _zz_338;
  wire                _zz_339;
  wire                _zz_340;
  wire                _zz_341;
  wire                _zz_342;
  wire                _zz_343;
  wire                _zz_344;
  wire                _zz_345;
  wire                _zz_346;
  wire                _zz_347;
  wire       [5:0]    _zz_cntLkHoldWrRmt_0_1;
  wire       [5:0]    _zz_cntLkHoldWrRmt_0_2;
  wire       [5:0]    _zz_cntLkWaitRmt_0_1;
  wire       [63:0]   _zz_348;
  wire       [5:0]    _zz_cntLkRespRmt_0_2;
  wire       [5:0]    _zz_cntRlseRespRmt_0_1;
  wire                when_TxnManCS_l303;
  wire                io_rdRmt_fire;
  wire                when_TxnManCS_l315;
  reg        [1:0]    compTxnCmtLoc_stateReg;
  reg        [1:0]    compTxnCmtLoc_stateNext;
  wire                when_TxnManCS_l369;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire       [5:0]    _zz_cntCmtReqLoc_0_1;
  reg        [1:0]    compLkRlseLoc_stateReg;
  reg        [1:0]    compLkRlseLoc_stateNext;
  wire       [5:0]    _zz_cntRlseReqWrLoc_0;
  wire       [63:0]   _zz_349;
  wire       [5:0]    _zz_when_TxnManCS_l440;
  wire                when_TxnManCS_l440;
  wire                lkReqRlseLoc_fire;
  wire       [5:0]    _zz_cntRlseReqLoc_0_1;
  wire                lkReqRlseLoc_fire_1;
  wire                when_TxnManCS_l456;
  wire       [5:0]    _zz_cntRlseReqWrLoc_0_1;
  reg        [1:0]    compLkRlseRmt_stateReg;
  reg        [1:0]    compLkRlseRmt_stateNext;
  wire       [5:0]    _zz_when_TxnManCS_l489;
  wire                when_TxnManCS_l489;
  wire                lkReqRlseRmt_fire;
  wire                when_TxnManCS_l505;
  wire       [63:0]   _zz_350;
  wire       [5:0]    _zz_cntRlseReqWrRmt_0;
  wire       [5:0]    _zz_cntRlseReqRmt_0_1;
  wire                io_wrRmt_fire;
  wire                when_TxnManCS_l521;
  wire       [5:0]    _zz_cntRlseReqRmt_0_2;
  reg        [1:0]    compTimeOut_stateReg;
  reg        [1:0]    compTimeOut_stateNext;
  wire                when_TxnManCS_l555;
  wire                when_TxnManCS_l555_1;
  wire                when_TxnManCS_l555_2;
  wire                when_TxnManCS_l555_3;
  wire                when_TxnManCS_l555_4;
  wire                when_TxnManCS_l555_5;
  wire                when_TxnManCS_l555_6;
  wire                when_TxnManCS_l555_7;
  wire                when_TxnManCS_l555_8;
  wire                when_TxnManCS_l555_9;
  wire                when_TxnManCS_l555_10;
  wire                when_TxnManCS_l555_11;
  wire                when_TxnManCS_l555_12;
  wire                when_TxnManCS_l555_13;
  wire                when_TxnManCS_l555_14;
  wire                when_TxnManCS_l555_15;
  wire                when_TxnManCS_l555_16;
  wire                when_TxnManCS_l555_17;
  wire                when_TxnManCS_l555_18;
  wire                when_TxnManCS_l555_19;
  wire                when_TxnManCS_l555_20;
  wire                when_TxnManCS_l555_21;
  wire                when_TxnManCS_l555_22;
  wire                when_TxnManCS_l555_23;
  wire                when_TxnManCS_l555_24;
  wire                when_TxnManCS_l555_25;
  wire                when_TxnManCS_l555_26;
  wire                when_TxnManCS_l555_27;
  wire                when_TxnManCS_l555_28;
  wire                when_TxnManCS_l555_29;
  wire                when_TxnManCS_l555_30;
  wire                when_TxnManCS_l555_31;
  wire                when_TxnManCS_l555_32;
  wire                when_TxnManCS_l555_33;
  wire                when_TxnManCS_l555_34;
  wire                when_TxnManCS_l555_35;
  wire                when_TxnManCS_l555_36;
  wire                when_TxnManCS_l555_37;
  wire                when_TxnManCS_l555_38;
  wire                when_TxnManCS_l555_39;
  wire                when_TxnManCS_l555_40;
  wire                when_TxnManCS_l555_41;
  wire                when_TxnManCS_l555_42;
  wire                when_TxnManCS_l555_43;
  wire                when_TxnManCS_l555_44;
  wire                when_TxnManCS_l555_45;
  wire                when_TxnManCS_l555_46;
  wire                when_TxnManCS_l555_47;
  wire                when_TxnManCS_l555_48;
  wire                when_TxnManCS_l555_49;
  wire                when_TxnManCS_l555_50;
  wire                when_TxnManCS_l555_51;
  wire                when_TxnManCS_l555_52;
  wire                when_TxnManCS_l555_53;
  wire                when_TxnManCS_l555_54;
  wire                when_TxnManCS_l555_55;
  wire                when_TxnManCS_l555_56;
  wire                when_TxnManCS_l555_57;
  wire                when_TxnManCS_l555_58;
  wire                when_TxnManCS_l555_59;
  wire                when_TxnManCS_l555_60;
  wire                when_TxnManCS_l555_61;
  wire                when_TxnManCS_l555_62;
  wire                when_TxnManCS_l555_63;
  reg        [2:0]    compLoadTxn_stateReg;
  reg        [2:0]    compLoadTxn_stateNext;
  wire                when_TxnManCS_l621;
  wire       [63:0]   _zz_351;
  wire                io_cmdAxi_ar_fire;
  wire                io_cmdAxi_r_fire_2;
  wire       [1:0]    _zz_352;
  wire       [1:0]    _zz_353;
  wire       [63:0]   _zz_354;
  wire       [63:0]   _zz_355;
  wire       [63:0]   _zz_356;
  wire       [63:0]   _zz_357;
  wire       [63:0]   _zz_358;
  wire       [63:0]   _zz_359;
  wire       [63:0]   _zz_360;
  wire       [63:0]   _zz_361;
  wire       [63:0]   _zz_362;
  wire       [63:0]   _zz_363;
  wire       [63:0]   _zz_364;
  wire       [63:0]   _zz_365;
  wire       [63:0]   _zz_366;
  wire       [63:0]   _zz_367;
  wire       [63:0]   _zz_368;
  wire       [63:0]   _zz_369;
  wire       [63:0]   _zz_370;
  wire       [63:0]   _zz_371;
  wire       [63:0]   _zz_372;
  wire       [63:0]   _zz_373;
  wire       [63:0]   _zz_374;
  wire       [63:0]   _zz_375;
  wire       [63:0]   _zz_376;
  wire       [63:0]   _zz_377;
  wire       [63:0]   _zz_378;
  wire       [63:0]   _zz_379;
  wire                when_TxnManCS_l665;
  reg        [1:0]    clkCnt_stateReg;
  reg        [1:0]    clkCnt_stateNext;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReqLoc_payload_lkType_string;
  reg [47:0] io_lkReqRmt_payload_lkType_string;
  reg [47:0] io_lkRespLoc_payload_lkType_string;
  reg [71:0] io_lkRespLoc_payload_respType_string;
  reg [47:0] io_lkRespRmt_payload_lkType_string;
  reg [71:0] io_lkRespRmt_payload_respType_string;
  reg [47:0] lkReqGetLoc_payload_lkType_string;
  reg [47:0] lkReqRlseLoc_payload_lkType_string;
  reg [47:0] lkReqGetRmt_payload_lkType_string;
  reg [47:0] lkReqRlseRmt_payload_lkType_string;
  reg [47:0] streamArbiter_8_io_output_s2mPipe_payload_lkType_string;
  reg [47:0] streamArbiter_8_io_output_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_string;
  reg [47:0] streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamArbiter_8_io_output_s2mPipe_rData_lkType_string;
  reg [47:0] streamArbiter_9_io_output_s2mPipe_payload_lkType_string;
  reg [47:0] streamArbiter_9_io_output_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_1_string;
  reg [47:0] streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamArbiter_9_io_output_s2mPipe_rData_lkType_string;
  reg [47:0] compLkReq_txnMemRd_payload_lkType_string;
  reg [47:0] _zz_compLkReq_txnMemRd_payload_lkType_string;
  reg [47:0] _zz_compLkReq_txnMemRd_payload_lkType_1_string;
  reg [47:0] _zz_lkReqGetLoc_payload_lkType_string;
  reg [47:0] _zz_lkReqGetRmt_payload_lkType_string;
  reg [47:0] compLkRespLoc_rLkResp_payload_lkType_string;
  reg [71:0] compLkRespLoc_rLkResp_payload_respType_string;
  reg [47:0] compLkRespRmt_rLkResp_payload_lkType_string;
  reg [71:0] compLkRespRmt_rLkResp_payload_respType_string;
  reg [47:0] compTxnCmtLoc_cmtTxn_lkType_string;
  reg [47:0] _zz_compTxnCmtLoc_cmtTxn_lkType_string;
  reg [47:0] compTxnCmtLoc_rCmtTxn_lkType_string;
  reg [47:0] compLkRlseLoc_lkItem_lkType_string;
  reg [71:0] compLkRlseLoc_lkItem_respType_string;
  reg [47:0] _zz_compLkRlseLoc_lkItem_lkType_string;
  reg [71:0] _zz_compLkRlseLoc_lkItem_respType_string;
  reg [47:0] _zz_lkReqRlseLoc_payload_lkType_string;
  reg [47:0] compLkRlseRmt_lkItem_lkType_string;
  reg [71:0] compLkRlseRmt_lkItem_respType_string;
  reg [47:0] _zz_compLkRlseRmt_lkItem_lkType_string;
  reg [71:0] _zz_compLkRlseRmt_lkItem_respType_string;
  reg [47:0] _zz_lkReqRlseRmt_payload_lkType_string;
  reg [47:0] compLkReq_stateReg_string;
  reg [47:0] compLkReq_stateNext_string;
  reg [95:0] compLkRespLoc_stateReg_string;
  reg [95:0] compLkRespLoc_stateNext_string;
  reg [111:0] compLkRespRmt_stateReg_string;
  reg [111:0] compLkRespRmt_stateNext_string;
  reg [63:0] compTxnCmtLoc_stateReg_string;
  reg [63:0] compTxnCmtLoc_stateNext_string;
  reg [55:0] compLkRlseLoc_stateReg_string;
  reg [55:0] compLkRlseLoc_stateNext_string;
  reg [87:0] compLkRlseRmt_stateReg_string;
  reg [87:0] compLkRlseRmt_stateNext_string;
  reg [39:0] compTimeOut_stateReg_string;
  reg [39:0] compTimeOut_stateNext_string;
  reg [71:0] compLoadTxn_stateReg_string;
  reg [71:0] compLoadTxn_stateNext_string;
  reg [47:0] _zz_352_string;
  reg [47:0] _zz_353_string;
  reg [31:0] clkCnt_stateReg_string;
  reg [31:0] clkCnt_stateNext_string;
  `endif

  reg [30:0] txnMem [0:4095];
  reg [30:0] txnWrMemLoc [0:4095];
  reg [30:0] txnWrMemRmt [0:4095];
  reg [48:0] lkMemLoc [0:4095];
  reg [48:0] lkMemRmt [0:4095];

  assign _zz_compLkReq_mskTxn2Start_ohFirst_masked = (compLkReq_mskTxn2Start_ohFirst_input - 64'h0000000000000001);
  assign _zz_compLkRespLoc_getAllRlseTimeOut = (_zz_cntLkHoldLoc_0 + _zz_cntLkWaitLoc_0);
  assign _zz_compLkRespLoc_getAllRlseTimeOut_2 = (_zz_compLkRespLoc_getAllRlseTimeOut_3 + _zz_compLkRespLoc_getAllRlseTimeOut_4);
  assign _zz_io_axi_ar_payload_addr = (_zz_io_axi_ar_payload_addr_1 + 28'h0);
  assign _zz_io_axi_ar_payload_addr_1 = ({6'd0,compLkRespLoc_rLkResp_payload_tId} <<< 6);
  assign _zz_io_axi_ar_payload_len = ({7'd0,1'b1} <<< compLkRespLoc_rLkResp_payload_wLen);
  assign _zz_compLkRespRmt_getAllRlseTimeOut_1 = (_zz_compLkRespRmt_getAllRlseTimeOut_2 + _zz_compLkRespRmt_getAllRlseTimeOut_3);
  assign _zz_compLkRespRmt_getAllRlseTimeOut_4 = (_zz_cntLkHoldRmt_0 + _zz_cntLkWaitRmt_0);
  assign _zz__zz_compTxnCmtLoc_cmtTxn_nId = {6'd0, _zz_cntCmtReqLoc_0};
  assign _zz_io_axi_aw_payload_addr = (_zz_io_axi_aw_payload_addr_1 + 28'h0);
  assign _zz_io_axi_aw_payload_addr_1 = ({6'd0,compTxnCmtLoc_cmtTxn_tId} <<< 6);
  assign _zz_io_axi_aw_payload_len = ({7'd0,1'b1} <<< compTxnCmtLoc_cmtTxn_wLen);
  assign _zz_io_axi_w_payload_last = (_zz_io_axi_w_payload_last_1 - 8'h01);
  assign _zz_io_axi_w_payload_last_1 = ({7'd0,1'b1} <<< compTxnCmtLoc_rCmtTxn_wLen);
  assign _zz__zz_compLkRlseLoc_lkItem_nId = {6'd0, _zz_cntRlseReqLoc_0};
  assign _zz__zz_compLkRlseRmt_lkItem_nId = {6'd0, _zz_cntRlseReqRmt_0};
  assign _zz_io_cmdAxi_ar_payload_addr = (_zz_io_cmdAxi_ar_payload_addr_1 + _zz_io_cmdAxi_ar_payload_addr_3);
  assign _zz_io_cmdAxi_ar_payload_addr_1 = ({3'd0,_zz_io_cmdAxi_ar_payload_addr_2} <<< 3);
  assign _zz_io_cmdAxi_ar_payload_addr_2 = ({6'd0,compLoadTxn_cntTxn} <<< 6);
  assign _zz_io_cmdAxi_ar_payload_addr_4 = ({6'd0,io_cmdAddrOffs} <<< 6);
  assign _zz_io_cmdAxi_ar_payload_addr_3 = {3'd0, _zz_io_cmdAxi_ar_payload_addr_4};
  assign _zz_io_cmdAxi_ar_payload_len = (_zz_io_cmdAxi_ar_payload_len_1 - 4'b0001);
  assign _zz_io_cmdAxi_ar_payload_len_1 = ({3'd0,1'b1} <<< 3);
  assign _zz_compLoadTxn_cntTxnWordInLine_valueNext_1 = compLoadTxn_cntTxnWordInLine_willIncrement;
  assign _zz_compLoadTxn_cntTxnWordInLine_valueNext = {2'd0, _zz_compLoadTxn_cntTxnWordInLine_valueNext_1};
  assign _zz_compLoadTxn_cntTxnWord_valueNext_1 = compLoadTxn_cntTxnWord_willIncrement;
  assign _zz_compLoadTxn_cntTxnWord_valueNext = {5'd0, _zz_compLoadTxn_cntTxnWord_valueNext_1};
  assign _zz_txnWrMemLoc_port_1 = (compLkReq_txnOffs + _zz_txnWrMemLoc_port_2);
  assign _zz_txnWrMemLoc_port_2 = {6'd0, _zz_cntLkReqWrLoc_0};
  assign _zz_txnWrMemRmt_port = (compLkReq_txnOffs + _zz_txnWrMemRmt_port_1);
  assign _zz_txnWrMemRmt_port_1 = {6'd0, _zz_cntLkReqWrRmt_0};
  assign _zz_compLkReq_txnLen = {compLkReq_txnMemRd_payload_wLen,{compLkReq_txnMemRd_payload_lkType,{compLkReq_txnMemRd_payload_tabId,{compLkReq_txnMemRd_payload_tId,compLkReq_txnMemRd_payload_nId}}}};
  assign _zz__zz_compLkReq_txnMemRdCmd_payload = (compLkReq_txnOffs + _zz__zz_compLkReq_txnMemRdCmd_payload_1);
  assign _zz__zz_compLkReq_txnMemRdCmd_payload_1 = {6'd0, compLkReq_reqIdx};
  assign _zz_compLkReq_txnMemRdCmd_payload_1 = (_zz_compLkReq_txnMemRdCmd_payload + 12'h001);
  assign _zz_when_TxnManCS_l128 = (compLkReq_txnLen - 6'h01);
  assign _zz_lkMemLoc_port_1 = (_zz_lkMemLoc_port_2 + _zz_lkMemLoc_port_4);
  assign _zz_lkMemLoc_port_2 = (compLkRespLoc_txnOffs + _zz_lkMemLoc_port_3);
  assign _zz_lkMemLoc_port_3 = {6'd0, _zz_cntLkHoldLoc_0};
  assign _zz_lkMemLoc_port_4 = {6'd0, _zz_cntLkWaitLoc_0};
  assign _zz_lkMemRmt_port_1 = (_zz_lkMemRmt_port_2 + _zz_lkMemRmt_port_4);
  assign _zz_lkMemRmt_port_2 = (compLkRespRmt_txnOffs + _zz_lkMemRmt_port_3);
  assign _zz_lkMemRmt_port_3 = {6'd0, _zz_cntLkHoldRmt_0};
  assign _zz_lkMemRmt_port_4 = {6'd0, _zz_cntLkWaitRmt_0};
  assign _zz_when_TxnManCS_l315 = (_zz_when_TxnManCS_l315_1 - 8'h01);
  assign _zz_when_TxnManCS_l315_1 = ({7'd0,1'b1} <<< compLkRespRmt_rLkResp_payload_wLen);
  assign _zz_when_TxnManCS_l440_3 = (_zz_when_TxnManCS_l440 + _zz_when_TxnManCS_l440_4);
  assign _zz_when_TxnManCS_l489_2 = (_zz_when_TxnManCS_l489 + _zz_when_TxnManCS_l489_3);
  assign _zz_when_TxnManCS_l521 = (_zz_when_TxnManCS_l521_1 - 8'h01);
  assign _zz_when_TxnManCS_l521_1 = ({7'd0,1'b1} <<< compLkRlseRmt_lkItem_wLen);
  assign _zz_txnMem_port = (compLoadTxn_txnOffs + _zz_txnMem_port_1);
  assign _zz_txnMem_port_1 = {6'd0, compLoadTxn_cntTxnWord_value};
  assign _zz_when_TxnManCS_l665 = (io_txnNumTotal - 32'h00000001);
  assign _zz_txnMem_port_2 = {compLoadTxn_txnBuff[30 : 28],{_zz_352,{compLoadTxn_txnBuff[25 : 23],{compLoadTxn_txnBuff[22 : 1],compLoadTxn_txnBuff[0 : 0]}}}};
  assign _zz__zz_compTxnCmtLoc_cmtTxn_nId_1 = 1'b1;
  assign _zz_txnWrMemLoc_port_3 = {compLkReq_txnMemRd_payload_wLen,{compLkReq_txnMemRd_payload_lkType,{compLkReq_txnMemRd_payload_tabId,{compLkReq_txnMemRd_payload_tId,compLkReq_txnMemRd_payload_nId}}}};
  assign _zz_txnWrMemRmt_port_2 = {compLkReq_txnMemRd_payload_wLen,{compLkReq_txnMemRd_payload_lkType,{compLkReq_txnMemRd_payload_tabId,{compLkReq_txnMemRd_payload_tId,compLkReq_txnMemRd_payload_nId}}}};
  assign _zz__zz_compLkRlseLoc_lkItem_nId_1 = 1'b1;
  assign _zz_lkMemLoc_port_5 = {io_lkRespLoc_payload_lkWaited,{io_lkRespLoc_payload_respType,{io_lkRespLoc_payload_wLen,{io_lkRespLoc_payload_lkIdx,{io_lkRespLoc_payload_txnAbt,{io_lkRespLoc_payload_lkRelease,{io_lkRespLoc_payload_lkType,{io_lkRespLoc_payload_txnId,{io_lkRespLoc_payload_snId,{io_lkRespLoc_payload_tabId,{io_lkRespLoc_payload_tId,io_lkRespLoc_payload_nId}}}}}}}}}}};
  assign _zz__zz_compLkRlseRmt_lkItem_nId_1 = 1'b1;
  assign _zz_lkMemRmt_port_5 = {io_lkRespRmt_payload_lkWaited,{io_lkRespRmt_payload_respType,{io_lkRespRmt_payload_wLen,{io_lkRespRmt_payload_lkIdx,{io_lkRespRmt_payload_txnAbt,{io_lkRespRmt_payload_lkRelease,{io_lkRespRmt_payload_lkType,{io_lkRespRmt_payload_txnId,{io_lkRespRmt_payload_snId,{io_lkRespRmt_payload_tabId,{io_lkRespRmt_payload_tId,io_lkRespRmt_payload_nId}}}}}}}}}}};
  assign _zz_compLkReq_mskTxn2Start = rReqDone_59;
  assign _zz_compLkReq_mskTxn2Start_1 = {rReqDone_58,{rReqDone_57,{rReqDone_56,{rReqDone_55,{rReqDone_54,{_zz_compLkReq_mskTxn2Start_2,_zz_compLkReq_mskTxn2Start_3}}}}}};
  assign _zz_compLkReq_mskTxn2Start_20 = rAbort_59;
  assign _zz_compLkReq_mskTxn2Start_21 = {rAbort_58,{rAbort_57,{rAbort_56,{rAbort_55,{rAbort_54,{_zz_compLkReq_mskTxn2Start_22,_zz_compLkReq_mskTxn2Start_23}}}}}};
  assign _zz_compLkReq_mskTxn2Start_2 = rReqDone_53;
  assign _zz_compLkReq_mskTxn2Start_3 = {rReqDone_52,{rReqDone_51,{rReqDone_50,{rReqDone_49,{rReqDone_48,{_zz_compLkReq_mskTxn2Start_4,_zz_compLkReq_mskTxn2Start_5}}}}}};
  assign _zz_compLkReq_mskTxn2Start_22 = rAbort_53;
  assign _zz_compLkReq_mskTxn2Start_23 = {rAbort_52,{rAbort_51,{rAbort_50,{rAbort_49,{rAbort_48,{_zz_compLkReq_mskTxn2Start_24,_zz_compLkReq_mskTxn2Start_25}}}}}};
  assign _zz_compLkReq_mskTxn2Start_4 = rReqDone_47;
  assign _zz_compLkReq_mskTxn2Start_5 = {rReqDone_46,{rReqDone_45,{rReqDone_44,{rReqDone_43,{rReqDone_42,{_zz_compLkReq_mskTxn2Start_6,_zz_compLkReq_mskTxn2Start_7}}}}}};
  assign _zz_compLkReq_mskTxn2Start_24 = rAbort_47;
  assign _zz_compLkReq_mskTxn2Start_25 = {rAbort_46,{rAbort_45,{rAbort_44,{rAbort_43,{rAbort_42,{_zz_compLkReq_mskTxn2Start_26,_zz_compLkReq_mskTxn2Start_27}}}}}};
  assign _zz_compLkReq_mskTxn2Start_6 = rReqDone_41;
  assign _zz_compLkReq_mskTxn2Start_7 = {rReqDone_40,{rReqDone_39,{rReqDone_38,{rReqDone_37,{rReqDone_36,{_zz_compLkReq_mskTxn2Start_8,_zz_compLkReq_mskTxn2Start_9}}}}}};
  assign _zz_compLkReq_mskTxn2Start_26 = rAbort_41;
  assign _zz_compLkReq_mskTxn2Start_27 = {rAbort_40,{rAbort_39,{rAbort_38,{rAbort_37,{rAbort_36,{_zz_compLkReq_mskTxn2Start_28,_zz_compLkReq_mskTxn2Start_29}}}}}};
  assign _zz_compLkReq_mskTxn2Start_8 = rReqDone_35;
  assign _zz_compLkReq_mskTxn2Start_9 = {rReqDone_34,{rReqDone_33,{rReqDone_32,{rReqDone_31,{rReqDone_30,{_zz_compLkReq_mskTxn2Start_10,_zz_compLkReq_mskTxn2Start_11}}}}}};
  assign _zz_compLkReq_mskTxn2Start_28 = rAbort_35;
  assign _zz_compLkReq_mskTxn2Start_29 = {rAbort_34,{rAbort_33,{rAbort_32,{rAbort_31,{rAbort_30,{_zz_compLkReq_mskTxn2Start_30,_zz_compLkReq_mskTxn2Start_31}}}}}};
  assign _zz_compLkReq_mskTxn2Start_10 = rReqDone_29;
  assign _zz_compLkReq_mskTxn2Start_11 = {rReqDone_28,{rReqDone_27,{rReqDone_26,{rReqDone_25,{rReqDone_24,{_zz_compLkReq_mskTxn2Start_12,_zz_compLkReq_mskTxn2Start_13}}}}}};
  assign _zz_compLkReq_mskTxn2Start_30 = rAbort_29;
  assign _zz_compLkReq_mskTxn2Start_31 = {rAbort_28,{rAbort_27,{rAbort_26,{rAbort_25,{rAbort_24,{_zz_compLkReq_mskTxn2Start_32,_zz_compLkReq_mskTxn2Start_33}}}}}};
  assign _zz_compLkReq_mskTxn2Start_12 = rReqDone_23;
  assign _zz_compLkReq_mskTxn2Start_13 = {rReqDone_22,{rReqDone_21,{rReqDone_20,{rReqDone_19,{rReqDone_18,{_zz_compLkReq_mskTxn2Start_14,_zz_compLkReq_mskTxn2Start_15}}}}}};
  assign _zz_compLkReq_mskTxn2Start_32 = rAbort_23;
  assign _zz_compLkReq_mskTxn2Start_33 = {rAbort_22,{rAbort_21,{rAbort_20,{rAbort_19,{rAbort_18,{_zz_compLkReq_mskTxn2Start_34,_zz_compLkReq_mskTxn2Start_35}}}}}};
  assign _zz_compLkReq_mskTxn2Start_14 = rReqDone_17;
  assign _zz_compLkReq_mskTxn2Start_15 = {rReqDone_16,{rReqDone_15,{rReqDone_14,{rReqDone_13,{rReqDone_12,{_zz_compLkReq_mskTxn2Start_16,_zz_compLkReq_mskTxn2Start_17}}}}}};
  assign _zz_compLkReq_mskTxn2Start_34 = rAbort_17;
  assign _zz_compLkReq_mskTxn2Start_35 = {rAbort_16,{rAbort_15,{rAbort_14,{rAbort_13,{rAbort_12,{_zz_compLkReq_mskTxn2Start_36,_zz_compLkReq_mskTxn2Start_37}}}}}};
  assign _zz_compLkReq_mskTxn2Start_16 = rReqDone_11;
  assign _zz_compLkReq_mskTxn2Start_17 = {rReqDone_10,{rReqDone_9,{rReqDone_8,{rReqDone_7,{rReqDone_6,{_zz_compLkReq_mskTxn2Start_18,_zz_compLkReq_mskTxn2Start_19}}}}}};
  assign _zz_compLkReq_mskTxn2Start_36 = rAbort_11;
  assign _zz_compLkReq_mskTxn2Start_37 = {rAbort_10,{rAbort_9,{rAbort_8,{rAbort_7,{rAbort_6,{_zz_compLkReq_mskTxn2Start_38,_zz_compLkReq_mskTxn2Start_39}}}}}};
  assign _zz_compLkReq_mskTxn2Start_18 = rReqDone_5;
  assign _zz_compLkReq_mskTxn2Start_19 = {rReqDone_4,{rReqDone_3,{rReqDone_2,{rReqDone_1,rReqDone_0}}}};
  assign _zz_compLkReq_mskTxn2Start_38 = rAbort_5;
  assign _zz_compLkReq_mskTxn2Start_39 = {rAbort_4,{rAbort_3,{rAbort_2,{rAbort_1,rAbort_0}}}};
  assign _zz__zz_compLkReq_rIdxTxn2Start_57 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[1] || _zz_compLkReq_rIdxTxn2Start) || _zz_compLkReq_rIdxTxn2Start_1) || _zz_compLkReq_rIdxTxn2Start_3) || _zz_compLkReq_rIdxTxn2Start_4) || _zz_compLkReq_rIdxTxn2Start_6) || _zz_compLkReq_rIdxTxn2Start_8) || _zz_compLkReq_rIdxTxn2Start_10) || _zz_compLkReq_rIdxTxn2Start_11) || _zz_compLkReq_rIdxTxn2Start_13) || _zz_compLkReq_rIdxTxn2Start_15) || _zz_compLkReq_rIdxTxn2Start_17) || _zz_compLkReq_rIdxTxn2Start_19) || _zz_compLkReq_rIdxTxn2Start_21) || _zz_compLkReq_rIdxTxn2Start_23) || _zz_compLkReq_rIdxTxn2Start_25);
  assign _zz__zz_compLkReq_rIdxTxn2Start_58 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[2] || _zz_compLkReq_rIdxTxn2Start) || _zz_compLkReq_rIdxTxn2Start_2) || _zz_compLkReq_rIdxTxn2Start_3) || _zz_compLkReq_rIdxTxn2Start_5) || _zz_compLkReq_rIdxTxn2Start_6) || _zz_compLkReq_rIdxTxn2Start_9) || _zz_compLkReq_rIdxTxn2Start_10) || _zz_compLkReq_rIdxTxn2Start_12) || _zz_compLkReq_rIdxTxn2Start_13) || _zz_compLkReq_rIdxTxn2Start_16) || _zz_compLkReq_rIdxTxn2Start_17) || _zz_compLkReq_rIdxTxn2Start_20) || _zz_compLkReq_rIdxTxn2Start_21) || _zz_compLkReq_rIdxTxn2Start_24) || _zz_compLkReq_rIdxTxn2Start_25);
  assign _zz__zz_compLkReq_rIdxTxn2Start_59 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[4] || _zz_compLkReq_rIdxTxn2Start_1) || _zz_compLkReq_rIdxTxn2Start_2) || _zz_compLkReq_rIdxTxn2Start_3) || _zz_compLkReq_rIdxTxn2Start_7) || _zz_compLkReq_rIdxTxn2Start_8) || _zz_compLkReq_rIdxTxn2Start_9) || _zz_compLkReq_rIdxTxn2Start_10) || _zz_compLkReq_rIdxTxn2Start_14) || _zz_compLkReq_rIdxTxn2Start_15) || _zz_compLkReq_rIdxTxn2Start_16) || _zz_compLkReq_rIdxTxn2Start_17) || _zz_compLkReq_rIdxTxn2Start_22) || _zz_compLkReq_rIdxTxn2Start_23) || _zz_compLkReq_rIdxTxn2Start_24) || _zz_compLkReq_rIdxTxn2Start_25);
  assign _zz__zz_compLkReq_rIdxTxn2Start_60 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[8] || _zz_compLkReq_rIdxTxn2Start_4) || _zz_compLkReq_rIdxTxn2Start_5) || _zz_compLkReq_rIdxTxn2Start_6) || _zz_compLkReq_rIdxTxn2Start_7) || _zz_compLkReq_rIdxTxn2Start_8) || _zz_compLkReq_rIdxTxn2Start_9) || _zz_compLkReq_rIdxTxn2Start_10) || _zz_compLkReq_rIdxTxn2Start_18) || _zz_compLkReq_rIdxTxn2Start_19) || _zz_compLkReq_rIdxTxn2Start_20) || _zz_compLkReq_rIdxTxn2Start_21) || _zz_compLkReq_rIdxTxn2Start_22) || _zz_compLkReq_rIdxTxn2Start_23) || _zz_compLkReq_rIdxTxn2Start_24) || _zz_compLkReq_rIdxTxn2Start_25);
  assign _zz__zz_compLkReq_rIdxTxn2Start_61 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[16] || _zz_compLkReq_rIdxTxn2Start_11) || _zz_compLkReq_rIdxTxn2Start_12) || _zz_compLkReq_rIdxTxn2Start_13) || _zz_compLkReq_rIdxTxn2Start_14) || _zz_compLkReq_rIdxTxn2Start_15) || _zz_compLkReq_rIdxTxn2Start_16) || _zz_compLkReq_rIdxTxn2Start_17) || _zz_compLkReq_rIdxTxn2Start_18) || _zz_compLkReq_rIdxTxn2Start_19) || _zz_compLkReq_rIdxTxn2Start_20) || _zz_compLkReq_rIdxTxn2Start_21) || _zz_compLkReq_rIdxTxn2Start_22) || _zz_compLkReq_rIdxTxn2Start_23) || _zz_compLkReq_rIdxTxn2Start_24) || _zz_compLkReq_rIdxTxn2Start_25);
  assign _zz__zz_compLkReq_rIdxTxn2Start_62 = (((((((((((((((compLkReq_mskTxn2Start_ohFirst_value[32] || _zz_compLkReq_rIdxTxn2Start_26) || _zz_compLkReq_rIdxTxn2Start_27) || _zz_compLkReq_rIdxTxn2Start_28) || _zz_compLkReq_rIdxTxn2Start_29) || _zz_compLkReq_rIdxTxn2Start_30) || _zz_compLkReq_rIdxTxn2Start_31) || _zz_compLkReq_rIdxTxn2Start_32) || _zz_compLkReq_rIdxTxn2Start_33) || _zz_compLkReq_rIdxTxn2Start_34) || _zz_compLkReq_rIdxTxn2Start_35) || _zz_compLkReq_rIdxTxn2Start_36) || _zz_compLkReq_rIdxTxn2Start_37) || _zz_compLkReq_rIdxTxn2Start_38) || _zz_compLkReq_rIdxTxn2Start_39) || _zz_compLkReq_rIdxTxn2Start_40);
  assign _zz_when_TxnManCS_l672 = ((((((((((((((((_zz_when_TxnManCS_l672_1 && rRlseDone_36) && rRlseDone_37) && rRlseDone_38) && rRlseDone_39) && rRlseDone_40) && rRlseDone_41) && rRlseDone_42) && rRlseDone_43) && rRlseDone_44) && rRlseDone_45) && rRlseDone_46) && rRlseDone_47) && rRlseDone_48) && rRlseDone_49) && rRlseDone_50) && rRlseDone_51);
  assign _zz_when_TxnManCS_l672_1 = ((((((((((((((((_zz_when_TxnManCS_l672_2 && rRlseDone_20) && rRlseDone_21) && rRlseDone_22) && rRlseDone_23) && rRlseDone_24) && rRlseDone_25) && rRlseDone_26) && rRlseDone_27) && rRlseDone_28) && rRlseDone_29) && rRlseDone_30) && rRlseDone_31) && rRlseDone_32) && rRlseDone_33) && rRlseDone_34) && rRlseDone_35);
  assign _zz_when_TxnManCS_l672_2 = ((((((((((((((((_zz_when_TxnManCS_l672_3 && rRlseDone_4) && rRlseDone_5) && rRlseDone_6) && rRlseDone_7) && rRlseDone_8) && rRlseDone_9) && rRlseDone_10) && rRlseDone_11) && rRlseDone_12) && rRlseDone_13) && rRlseDone_14) && rRlseDone_15) && rRlseDone_16) && rRlseDone_17) && rRlseDone_18) && rRlseDone_19);
  assign _zz_when_TxnManCS_l672_3 = (((rRlseDone_0 && rRlseDone_1) && rRlseDone_2) && rRlseDone_3);
  always @(posedge clk) begin
    if(compLkReq_txnMemRdCmd_ready) begin
      _zz_txnMem_port0 <= txnMem[compLkReq_txnMemRdCmd_payload];
    end
  end

  always @(posedge clk) begin
    if(compLoadTxn_rTxnMemLd) begin
      txnMem[_zz_txnMem_port] <= _zz_txnMem_port_2;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_compTxnCmtLoc_cmtTxn_nId_1) begin
      _zz_txnWrMemLoc_port0 <= txnWrMemLoc[_zz_compTxnCmtLoc_cmtTxn_nId];
    end
  end

  always @(posedge clk) begin
    if(_zz_4) begin
      txnWrMemLoc[_zz_txnWrMemLoc_port_1] <= _zz_txnWrMemLoc_port_3;
    end
  end

  always @(posedge clk) begin
    if(_zz_3) begin
      txnWrMemRmt[_zz_txnWrMemRmt_port] <= _zz_txnWrMemRmt_port_2;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_compLkRlseLoc_lkItem_nId_1) begin
      _zz_lkMemLoc_port0 <= lkMemLoc[_zz_compLkRlseLoc_lkItem_nId];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      lkMemLoc[_zz_lkMemLoc_port_1] <= _zz_lkMemLoc_port_5;
    end
  end

  always @(posedge clk) begin
    if(_zz__zz_compLkRlseRmt_lkItem_nId_1) begin
      _zz_lkMemRmt_port0 <= lkMemRmt[_zz_compLkRlseRmt_lkItem_nId];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      lkMemRmt[_zz_lkMemRmt_port_1] <= _zz_lkMemRmt_port_5;
    end
  end

  StreamArbiter_5 streamArbiter_8 (
    .io_inputs_0_valid              (lkReqGetLoc_valid                            ), //i
    .io_inputs_0_ready              (streamArbiter_8_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_nId        (lkReqGetLoc_payload_nId                      ), //i
    .io_inputs_0_payload_tId        (lkReqGetLoc_payload_tId[21:0]                ), //i
    .io_inputs_0_payload_tabId      (lkReqGetLoc_payload_tabId[2:0]               ), //i
    .io_inputs_0_payload_snId       (lkReqGetLoc_payload_snId                     ), //i
    .io_inputs_0_payload_txnId      (lkReqGetLoc_payload_txnId[5:0]               ), //i
    .io_inputs_0_payload_lkType     (lkReqGetLoc_payload_lkType[1:0]              ), //i
    .io_inputs_0_payload_lkRelease  (lkReqGetLoc_payload_lkRelease                ), //i
    .io_inputs_0_payload_txnTimeOut (lkReqGetLoc_payload_txnTimeOut               ), //i
    .io_inputs_0_payload_txnAbt     (lkReqGetLoc_payload_txnAbt                   ), //i
    .io_inputs_0_payload_lkIdx      (lkReqGetLoc_payload_lkIdx[5:0]               ), //i
    .io_inputs_0_payload_wLen       (lkReqGetLoc_payload_wLen[2:0]                ), //i
    .io_inputs_1_valid              (lkReqRlseLoc_valid                           ), //i
    .io_inputs_1_ready              (streamArbiter_8_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_nId        (lkReqRlseLoc_payload_nId                     ), //i
    .io_inputs_1_payload_tId        (lkReqRlseLoc_payload_tId[21:0]               ), //i
    .io_inputs_1_payload_tabId      (lkReqRlseLoc_payload_tabId[2:0]              ), //i
    .io_inputs_1_payload_snId       (lkReqRlseLoc_payload_snId                    ), //i
    .io_inputs_1_payload_txnId      (lkReqRlseLoc_payload_txnId[5:0]              ), //i
    .io_inputs_1_payload_lkType     (lkReqRlseLoc_payload_lkType[1:0]             ), //i
    .io_inputs_1_payload_lkRelease  (lkReqRlseLoc_payload_lkRelease               ), //i
    .io_inputs_1_payload_txnTimeOut (lkReqRlseLoc_payload_txnTimeOut              ), //i
    .io_inputs_1_payload_txnAbt     (lkReqRlseLoc_payload_txnAbt                  ), //i
    .io_inputs_1_payload_lkIdx      (lkReqRlseLoc_payload_lkIdx[5:0]              ), //i
    .io_inputs_1_payload_wLen       (lkReqRlseLoc_payload_wLen[2:0]               ), //i
    .io_output_valid                (streamArbiter_8_io_output_valid              ), //o
    .io_output_ready                (streamArbiter_8_io_output_ready              ), //i
    .io_output_payload_nId          (streamArbiter_8_io_output_payload_nId        ), //o
    .io_output_payload_tId          (streamArbiter_8_io_output_payload_tId[21:0]  ), //o
    .io_output_payload_tabId        (streamArbiter_8_io_output_payload_tabId[2:0] ), //o
    .io_output_payload_snId         (streamArbiter_8_io_output_payload_snId       ), //o
    .io_output_payload_txnId        (streamArbiter_8_io_output_payload_txnId[5:0] ), //o
    .io_output_payload_lkType       (streamArbiter_8_io_output_payload_lkType[1:0]), //o
    .io_output_payload_lkRelease    (streamArbiter_8_io_output_payload_lkRelease  ), //o
    .io_output_payload_txnTimeOut   (streamArbiter_8_io_output_payload_txnTimeOut ), //o
    .io_output_payload_txnAbt       (streamArbiter_8_io_output_payload_txnAbt     ), //o
    .io_output_payload_lkIdx        (streamArbiter_8_io_output_payload_lkIdx[5:0] ), //o
    .io_output_payload_wLen         (streamArbiter_8_io_output_payload_wLen[2:0]  ), //o
    .io_chosen                      (streamArbiter_8_io_chosen                    ), //o
    .io_chosenOH                    (streamArbiter_8_io_chosenOH[1:0]             ), //o
    .clk                            (clk                                          ), //i
    .resetn                         (resetn                                       )  //i
  );
  StreamArbiter_5 streamArbiter_9 (
    .io_inputs_0_valid              (lkReqGetRmt_valid                            ), //i
    .io_inputs_0_ready              (streamArbiter_9_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_nId        (lkReqGetRmt_payload_nId                      ), //i
    .io_inputs_0_payload_tId        (lkReqGetRmt_payload_tId[21:0]                ), //i
    .io_inputs_0_payload_tabId      (lkReqGetRmt_payload_tabId[2:0]               ), //i
    .io_inputs_0_payload_snId       (lkReqGetRmt_payload_snId                     ), //i
    .io_inputs_0_payload_txnId      (lkReqGetRmt_payload_txnId[5:0]               ), //i
    .io_inputs_0_payload_lkType     (lkReqGetRmt_payload_lkType[1:0]              ), //i
    .io_inputs_0_payload_lkRelease  (lkReqGetRmt_payload_lkRelease                ), //i
    .io_inputs_0_payload_txnTimeOut (lkReqGetRmt_payload_txnTimeOut               ), //i
    .io_inputs_0_payload_txnAbt     (lkReqGetRmt_payload_txnAbt                   ), //i
    .io_inputs_0_payload_lkIdx      (lkReqGetRmt_payload_lkIdx[5:0]               ), //i
    .io_inputs_0_payload_wLen       (lkReqGetRmt_payload_wLen[2:0]                ), //i
    .io_inputs_1_valid              (lkReqRlseRmt_valid                           ), //i
    .io_inputs_1_ready              (streamArbiter_9_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_nId        (lkReqRlseRmt_payload_nId                     ), //i
    .io_inputs_1_payload_tId        (lkReqRlseRmt_payload_tId[21:0]               ), //i
    .io_inputs_1_payload_tabId      (lkReqRlseRmt_payload_tabId[2:0]              ), //i
    .io_inputs_1_payload_snId       (lkReqRlseRmt_payload_snId                    ), //i
    .io_inputs_1_payload_txnId      (lkReqRlseRmt_payload_txnId[5:0]              ), //i
    .io_inputs_1_payload_lkType     (lkReqRlseRmt_payload_lkType[1:0]             ), //i
    .io_inputs_1_payload_lkRelease  (lkReqRlseRmt_payload_lkRelease               ), //i
    .io_inputs_1_payload_txnTimeOut (lkReqRlseRmt_payload_txnTimeOut              ), //i
    .io_inputs_1_payload_txnAbt     (lkReqRlseRmt_payload_txnAbt                  ), //i
    .io_inputs_1_payload_lkIdx      (lkReqRlseRmt_payload_lkIdx[5:0]              ), //i
    .io_inputs_1_payload_wLen       (lkReqRlseRmt_payload_wLen[2:0]               ), //i
    .io_output_valid                (streamArbiter_9_io_output_valid              ), //o
    .io_output_ready                (streamArbiter_9_io_output_ready              ), //i
    .io_output_payload_nId          (streamArbiter_9_io_output_payload_nId        ), //o
    .io_output_payload_tId          (streamArbiter_9_io_output_payload_tId[21:0]  ), //o
    .io_output_payload_tabId        (streamArbiter_9_io_output_payload_tabId[2:0] ), //o
    .io_output_payload_snId         (streamArbiter_9_io_output_payload_snId       ), //o
    .io_output_payload_txnId        (streamArbiter_9_io_output_payload_txnId[5:0] ), //o
    .io_output_payload_lkType       (streamArbiter_9_io_output_payload_lkType[1:0]), //o
    .io_output_payload_lkRelease    (streamArbiter_9_io_output_payload_lkRelease  ), //o
    .io_output_payload_txnTimeOut   (streamArbiter_9_io_output_payload_txnTimeOut ), //o
    .io_output_payload_txnAbt       (streamArbiter_9_io_output_payload_txnAbt     ), //o
    .io_output_payload_lkIdx        (streamArbiter_9_io_output_payload_lkIdx[5:0] ), //o
    .io_output_payload_wLen         (streamArbiter_9_io_output_payload_wLen[2:0]  ), //o
    .io_chosen                      (streamArbiter_9_io_chosen                    ), //o
    .io_chosenOH                    (streamArbiter_9_io_chosenOH[1:0]             ), //o
    .clk                            (clk                                          ), //i
    .resetn                         (resetn                                       )  //i
  );
  always @(*) begin
    case(compLkRespLoc_rCurTxnId)
      6'b000000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_0;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_0;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_0;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_0;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_0;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_0;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_0;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_0;
        _zz_when_TxnManCS_l166 = rAbort_0;
        _zz_when_TxnManCS_l164 = rTimeOut_0;
        _zz_when_TxnManCS_l164_1 = rReqDone_0;
      end
      6'b000001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_1;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_1;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_1;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_1;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_1;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_1;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_1;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_1;
        _zz_when_TxnManCS_l166 = rAbort_1;
        _zz_when_TxnManCS_l164 = rTimeOut_1;
        _zz_when_TxnManCS_l164_1 = rReqDone_1;
      end
      6'b000010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_2;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_2;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_2;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_2;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_2;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_2;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_2;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_2;
        _zz_when_TxnManCS_l166 = rAbort_2;
        _zz_when_TxnManCS_l164 = rTimeOut_2;
        _zz_when_TxnManCS_l164_1 = rReqDone_2;
      end
      6'b000011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_3;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_3;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_3;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_3;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_3;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_3;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_3;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_3;
        _zz_when_TxnManCS_l166 = rAbort_3;
        _zz_when_TxnManCS_l164 = rTimeOut_3;
        _zz_when_TxnManCS_l164_1 = rReqDone_3;
      end
      6'b000100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_4;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_4;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_4;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_4;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_4;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_4;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_4;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_4;
        _zz_when_TxnManCS_l166 = rAbort_4;
        _zz_when_TxnManCS_l164 = rTimeOut_4;
        _zz_when_TxnManCS_l164_1 = rReqDone_4;
      end
      6'b000101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_5;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_5;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_5;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_5;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_5;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_5;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_5;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_5;
        _zz_when_TxnManCS_l166 = rAbort_5;
        _zz_when_TxnManCS_l164 = rTimeOut_5;
        _zz_when_TxnManCS_l164_1 = rReqDone_5;
      end
      6'b000110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_6;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_6;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_6;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_6;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_6;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_6;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_6;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_6;
        _zz_when_TxnManCS_l166 = rAbort_6;
        _zz_when_TxnManCS_l164 = rTimeOut_6;
        _zz_when_TxnManCS_l164_1 = rReqDone_6;
      end
      6'b000111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_7;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_7;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_7;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_7;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_7;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_7;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_7;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_7;
        _zz_when_TxnManCS_l166 = rAbort_7;
        _zz_when_TxnManCS_l164 = rTimeOut_7;
        _zz_when_TxnManCS_l164_1 = rReqDone_7;
      end
      6'b001000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_8;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_8;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_8;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_8;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_8;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_8;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_8;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_8;
        _zz_when_TxnManCS_l166 = rAbort_8;
        _zz_when_TxnManCS_l164 = rTimeOut_8;
        _zz_when_TxnManCS_l164_1 = rReqDone_8;
      end
      6'b001001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_9;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_9;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_9;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_9;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_9;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_9;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_9;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_9;
        _zz_when_TxnManCS_l166 = rAbort_9;
        _zz_when_TxnManCS_l164 = rTimeOut_9;
        _zz_when_TxnManCS_l164_1 = rReqDone_9;
      end
      6'b001010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_10;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_10;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_10;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_10;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_10;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_10;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_10;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_10;
        _zz_when_TxnManCS_l166 = rAbort_10;
        _zz_when_TxnManCS_l164 = rTimeOut_10;
        _zz_when_TxnManCS_l164_1 = rReqDone_10;
      end
      6'b001011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_11;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_11;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_11;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_11;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_11;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_11;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_11;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_11;
        _zz_when_TxnManCS_l166 = rAbort_11;
        _zz_when_TxnManCS_l164 = rTimeOut_11;
        _zz_when_TxnManCS_l164_1 = rReqDone_11;
      end
      6'b001100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_12;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_12;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_12;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_12;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_12;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_12;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_12;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_12;
        _zz_when_TxnManCS_l166 = rAbort_12;
        _zz_when_TxnManCS_l164 = rTimeOut_12;
        _zz_when_TxnManCS_l164_1 = rReqDone_12;
      end
      6'b001101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_13;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_13;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_13;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_13;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_13;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_13;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_13;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_13;
        _zz_when_TxnManCS_l166 = rAbort_13;
        _zz_when_TxnManCS_l164 = rTimeOut_13;
        _zz_when_TxnManCS_l164_1 = rReqDone_13;
      end
      6'b001110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_14;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_14;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_14;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_14;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_14;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_14;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_14;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_14;
        _zz_when_TxnManCS_l166 = rAbort_14;
        _zz_when_TxnManCS_l164 = rTimeOut_14;
        _zz_when_TxnManCS_l164_1 = rReqDone_14;
      end
      6'b001111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_15;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_15;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_15;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_15;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_15;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_15;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_15;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_15;
        _zz_when_TxnManCS_l166 = rAbort_15;
        _zz_when_TxnManCS_l164 = rTimeOut_15;
        _zz_when_TxnManCS_l164_1 = rReqDone_15;
      end
      6'b010000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_16;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_16;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_16;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_16;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_16;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_16;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_16;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_16;
        _zz_when_TxnManCS_l166 = rAbort_16;
        _zz_when_TxnManCS_l164 = rTimeOut_16;
        _zz_when_TxnManCS_l164_1 = rReqDone_16;
      end
      6'b010001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_17;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_17;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_17;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_17;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_17;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_17;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_17;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_17;
        _zz_when_TxnManCS_l166 = rAbort_17;
        _zz_when_TxnManCS_l164 = rTimeOut_17;
        _zz_when_TxnManCS_l164_1 = rReqDone_17;
      end
      6'b010010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_18;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_18;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_18;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_18;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_18;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_18;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_18;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_18;
        _zz_when_TxnManCS_l166 = rAbort_18;
        _zz_when_TxnManCS_l164 = rTimeOut_18;
        _zz_when_TxnManCS_l164_1 = rReqDone_18;
      end
      6'b010011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_19;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_19;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_19;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_19;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_19;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_19;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_19;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_19;
        _zz_when_TxnManCS_l166 = rAbort_19;
        _zz_when_TxnManCS_l164 = rTimeOut_19;
        _zz_when_TxnManCS_l164_1 = rReqDone_19;
      end
      6'b010100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_20;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_20;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_20;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_20;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_20;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_20;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_20;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_20;
        _zz_when_TxnManCS_l166 = rAbort_20;
        _zz_when_TxnManCS_l164 = rTimeOut_20;
        _zz_when_TxnManCS_l164_1 = rReqDone_20;
      end
      6'b010101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_21;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_21;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_21;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_21;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_21;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_21;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_21;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_21;
        _zz_when_TxnManCS_l166 = rAbort_21;
        _zz_when_TxnManCS_l164 = rTimeOut_21;
        _zz_when_TxnManCS_l164_1 = rReqDone_21;
      end
      6'b010110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_22;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_22;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_22;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_22;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_22;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_22;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_22;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_22;
        _zz_when_TxnManCS_l166 = rAbort_22;
        _zz_when_TxnManCS_l164 = rTimeOut_22;
        _zz_when_TxnManCS_l164_1 = rReqDone_22;
      end
      6'b010111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_23;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_23;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_23;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_23;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_23;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_23;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_23;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_23;
        _zz_when_TxnManCS_l166 = rAbort_23;
        _zz_when_TxnManCS_l164 = rTimeOut_23;
        _zz_when_TxnManCS_l164_1 = rReqDone_23;
      end
      6'b011000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_24;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_24;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_24;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_24;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_24;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_24;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_24;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_24;
        _zz_when_TxnManCS_l166 = rAbort_24;
        _zz_when_TxnManCS_l164 = rTimeOut_24;
        _zz_when_TxnManCS_l164_1 = rReqDone_24;
      end
      6'b011001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_25;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_25;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_25;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_25;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_25;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_25;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_25;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_25;
        _zz_when_TxnManCS_l166 = rAbort_25;
        _zz_when_TxnManCS_l164 = rTimeOut_25;
        _zz_when_TxnManCS_l164_1 = rReqDone_25;
      end
      6'b011010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_26;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_26;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_26;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_26;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_26;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_26;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_26;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_26;
        _zz_when_TxnManCS_l166 = rAbort_26;
        _zz_when_TxnManCS_l164 = rTimeOut_26;
        _zz_when_TxnManCS_l164_1 = rReqDone_26;
      end
      6'b011011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_27;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_27;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_27;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_27;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_27;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_27;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_27;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_27;
        _zz_when_TxnManCS_l166 = rAbort_27;
        _zz_when_TxnManCS_l164 = rTimeOut_27;
        _zz_when_TxnManCS_l164_1 = rReqDone_27;
      end
      6'b011100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_28;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_28;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_28;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_28;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_28;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_28;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_28;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_28;
        _zz_when_TxnManCS_l166 = rAbort_28;
        _zz_when_TxnManCS_l164 = rTimeOut_28;
        _zz_when_TxnManCS_l164_1 = rReqDone_28;
      end
      6'b011101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_29;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_29;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_29;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_29;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_29;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_29;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_29;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_29;
        _zz_when_TxnManCS_l166 = rAbort_29;
        _zz_when_TxnManCS_l164 = rTimeOut_29;
        _zz_when_TxnManCS_l164_1 = rReqDone_29;
      end
      6'b011110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_30;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_30;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_30;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_30;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_30;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_30;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_30;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_30;
        _zz_when_TxnManCS_l166 = rAbort_30;
        _zz_when_TxnManCS_l164 = rTimeOut_30;
        _zz_when_TxnManCS_l164_1 = rReqDone_30;
      end
      6'b011111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_31;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_31;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_31;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_31;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_31;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_31;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_31;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_31;
        _zz_when_TxnManCS_l166 = rAbort_31;
        _zz_when_TxnManCS_l164 = rTimeOut_31;
        _zz_when_TxnManCS_l164_1 = rReqDone_31;
      end
      6'b100000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_32;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_32;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_32;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_32;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_32;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_32;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_32;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_32;
        _zz_when_TxnManCS_l166 = rAbort_32;
        _zz_when_TxnManCS_l164 = rTimeOut_32;
        _zz_when_TxnManCS_l164_1 = rReqDone_32;
      end
      6'b100001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_33;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_33;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_33;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_33;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_33;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_33;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_33;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_33;
        _zz_when_TxnManCS_l166 = rAbort_33;
        _zz_when_TxnManCS_l164 = rTimeOut_33;
        _zz_when_TxnManCS_l164_1 = rReqDone_33;
      end
      6'b100010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_34;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_34;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_34;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_34;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_34;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_34;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_34;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_34;
        _zz_when_TxnManCS_l166 = rAbort_34;
        _zz_when_TxnManCS_l164 = rTimeOut_34;
        _zz_when_TxnManCS_l164_1 = rReqDone_34;
      end
      6'b100011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_35;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_35;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_35;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_35;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_35;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_35;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_35;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_35;
        _zz_when_TxnManCS_l166 = rAbort_35;
        _zz_when_TxnManCS_l164 = rTimeOut_35;
        _zz_when_TxnManCS_l164_1 = rReqDone_35;
      end
      6'b100100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_36;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_36;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_36;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_36;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_36;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_36;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_36;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_36;
        _zz_when_TxnManCS_l166 = rAbort_36;
        _zz_when_TxnManCS_l164 = rTimeOut_36;
        _zz_when_TxnManCS_l164_1 = rReqDone_36;
      end
      6'b100101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_37;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_37;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_37;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_37;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_37;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_37;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_37;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_37;
        _zz_when_TxnManCS_l166 = rAbort_37;
        _zz_when_TxnManCS_l164 = rTimeOut_37;
        _zz_when_TxnManCS_l164_1 = rReqDone_37;
      end
      6'b100110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_38;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_38;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_38;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_38;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_38;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_38;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_38;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_38;
        _zz_when_TxnManCS_l166 = rAbort_38;
        _zz_when_TxnManCS_l164 = rTimeOut_38;
        _zz_when_TxnManCS_l164_1 = rReqDone_38;
      end
      6'b100111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_39;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_39;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_39;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_39;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_39;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_39;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_39;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_39;
        _zz_when_TxnManCS_l166 = rAbort_39;
        _zz_when_TxnManCS_l164 = rTimeOut_39;
        _zz_when_TxnManCS_l164_1 = rReqDone_39;
      end
      6'b101000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_40;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_40;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_40;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_40;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_40;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_40;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_40;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_40;
        _zz_when_TxnManCS_l166 = rAbort_40;
        _zz_when_TxnManCS_l164 = rTimeOut_40;
        _zz_when_TxnManCS_l164_1 = rReqDone_40;
      end
      6'b101001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_41;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_41;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_41;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_41;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_41;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_41;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_41;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_41;
        _zz_when_TxnManCS_l166 = rAbort_41;
        _zz_when_TxnManCS_l164 = rTimeOut_41;
        _zz_when_TxnManCS_l164_1 = rReqDone_41;
      end
      6'b101010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_42;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_42;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_42;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_42;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_42;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_42;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_42;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_42;
        _zz_when_TxnManCS_l166 = rAbort_42;
        _zz_when_TxnManCS_l164 = rTimeOut_42;
        _zz_when_TxnManCS_l164_1 = rReqDone_42;
      end
      6'b101011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_43;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_43;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_43;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_43;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_43;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_43;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_43;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_43;
        _zz_when_TxnManCS_l166 = rAbort_43;
        _zz_when_TxnManCS_l164 = rTimeOut_43;
        _zz_when_TxnManCS_l164_1 = rReqDone_43;
      end
      6'b101100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_44;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_44;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_44;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_44;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_44;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_44;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_44;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_44;
        _zz_when_TxnManCS_l166 = rAbort_44;
        _zz_when_TxnManCS_l164 = rTimeOut_44;
        _zz_when_TxnManCS_l164_1 = rReqDone_44;
      end
      6'b101101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_45;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_45;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_45;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_45;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_45;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_45;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_45;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_45;
        _zz_when_TxnManCS_l166 = rAbort_45;
        _zz_when_TxnManCS_l164 = rTimeOut_45;
        _zz_when_TxnManCS_l164_1 = rReqDone_45;
      end
      6'b101110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_46;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_46;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_46;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_46;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_46;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_46;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_46;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_46;
        _zz_when_TxnManCS_l166 = rAbort_46;
        _zz_when_TxnManCS_l164 = rTimeOut_46;
        _zz_when_TxnManCS_l164_1 = rReqDone_46;
      end
      6'b101111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_47;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_47;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_47;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_47;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_47;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_47;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_47;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_47;
        _zz_when_TxnManCS_l166 = rAbort_47;
        _zz_when_TxnManCS_l164 = rTimeOut_47;
        _zz_when_TxnManCS_l164_1 = rReqDone_47;
      end
      6'b110000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_48;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_48;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_48;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_48;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_48;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_48;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_48;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_48;
        _zz_when_TxnManCS_l166 = rAbort_48;
        _zz_when_TxnManCS_l164 = rTimeOut_48;
        _zz_when_TxnManCS_l164_1 = rReqDone_48;
      end
      6'b110001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_49;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_49;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_49;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_49;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_49;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_49;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_49;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_49;
        _zz_when_TxnManCS_l166 = rAbort_49;
        _zz_when_TxnManCS_l164 = rTimeOut_49;
        _zz_when_TxnManCS_l164_1 = rReqDone_49;
      end
      6'b110010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_50;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_50;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_50;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_50;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_50;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_50;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_50;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_50;
        _zz_when_TxnManCS_l166 = rAbort_50;
        _zz_when_TxnManCS_l164 = rTimeOut_50;
        _zz_when_TxnManCS_l164_1 = rReqDone_50;
      end
      6'b110011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_51;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_51;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_51;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_51;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_51;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_51;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_51;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_51;
        _zz_when_TxnManCS_l166 = rAbort_51;
        _zz_when_TxnManCS_l164 = rTimeOut_51;
        _zz_when_TxnManCS_l164_1 = rReqDone_51;
      end
      6'b110100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_52;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_52;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_52;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_52;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_52;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_52;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_52;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_52;
        _zz_when_TxnManCS_l166 = rAbort_52;
        _zz_when_TxnManCS_l164 = rTimeOut_52;
        _zz_when_TxnManCS_l164_1 = rReqDone_52;
      end
      6'b110101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_53;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_53;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_53;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_53;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_53;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_53;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_53;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_53;
        _zz_when_TxnManCS_l166 = rAbort_53;
        _zz_when_TxnManCS_l164 = rTimeOut_53;
        _zz_when_TxnManCS_l164_1 = rReqDone_53;
      end
      6'b110110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_54;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_54;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_54;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_54;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_54;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_54;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_54;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_54;
        _zz_when_TxnManCS_l166 = rAbort_54;
        _zz_when_TxnManCS_l164 = rTimeOut_54;
        _zz_when_TxnManCS_l164_1 = rReqDone_54;
      end
      6'b110111 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_55;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_55;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_55;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_55;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_55;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_55;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_55;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_55;
        _zz_when_TxnManCS_l166 = rAbort_55;
        _zz_when_TxnManCS_l164 = rTimeOut_55;
        _zz_when_TxnManCS_l164_1 = rReqDone_55;
      end
      6'b111000 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_56;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_56;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_56;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_56;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_56;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_56;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_56;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_56;
        _zz_when_TxnManCS_l166 = rAbort_56;
        _zz_when_TxnManCS_l164 = rTimeOut_56;
        _zz_when_TxnManCS_l164_1 = rReqDone_56;
      end
      6'b111001 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_57;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_57;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_57;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_57;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_57;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_57;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_57;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_57;
        _zz_when_TxnManCS_l166 = rAbort_57;
        _zz_when_TxnManCS_l164 = rTimeOut_57;
        _zz_when_TxnManCS_l164_1 = rReqDone_57;
      end
      6'b111010 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_58;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_58;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_58;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_58;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_58;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_58;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_58;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_58;
        _zz_when_TxnManCS_l166 = rAbort_58;
        _zz_when_TxnManCS_l164 = rTimeOut_58;
        _zz_when_TxnManCS_l164_1 = rReqDone_58;
      end
      6'b111011 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_59;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_59;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_59;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_59;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_59;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_59;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_59;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_59;
        _zz_when_TxnManCS_l166 = rAbort_59;
        _zz_when_TxnManCS_l164 = rTimeOut_59;
        _zz_when_TxnManCS_l164_1 = rReqDone_59;
      end
      6'b111100 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_60;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_60;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_60;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_60;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_60;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_60;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_60;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_60;
        _zz_when_TxnManCS_l166 = rAbort_60;
        _zz_when_TxnManCS_l164 = rTimeOut_60;
        _zz_when_TxnManCS_l164_1 = rReqDone_60;
      end
      6'b111101 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_61;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_61;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_61;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_61;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_61;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_61;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_61;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_61;
        _zz_when_TxnManCS_l166 = rAbort_61;
        _zz_when_TxnManCS_l164 = rTimeOut_61;
        _zz_when_TxnManCS_l164_1 = rReqDone_61;
      end
      6'b111110 : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_62;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_62;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_62;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_62;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_62;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_62;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_62;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_62;
        _zz_when_TxnManCS_l166 = rAbort_62;
        _zz_when_TxnManCS_l164 = rTimeOut_62;
        _zz_when_TxnManCS_l164_1 = rReqDone_62;
      end
      default : begin
        _zz_compLkRespLoc_getAllRlse = cntRlseRespLoc_63;
        _zz_compLkRespLoc_getAllRlse_1 = cntLkHoldLoc_63;
        _zz_compLkRespLoc_getAllRlse_2 = cntRlseRespRmt_63;
        _zz_compLkRespLoc_getAllRlse_3 = cntLkHoldRmt_63;
        _zz_compLkRespLoc_getAllLkResp = cntLkReqLoc_63;
        _zz_compLkRespLoc_getAllLkResp_1 = cntLkRespLoc_63;
        _zz_compLkRespLoc_getAllLkResp_2 = cntLkReqRmt_63;
        _zz_compLkRespLoc_getAllLkResp_3 = cntLkRespRmt_63;
        _zz_when_TxnManCS_l166 = rAbort_63;
        _zz_when_TxnManCS_l164 = rTimeOut_63;
        _zz_when_TxnManCS_l164_1 = rReqDone_63;
      end
    endcase
  end

  always @(*) begin
    case(io_lkRespLoc_payload_txnId)
      6'b000000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_0;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_0;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_0;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_0;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_0;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_0;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_0;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_0;
      end
      6'b000001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_1;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_1;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_1;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_1;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_1;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_1;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_1;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_1;
      end
      6'b000010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_2;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_2;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_2;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_2;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_2;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_2;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_2;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_2;
      end
      6'b000011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_3;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_3;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_3;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_3;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_3;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_3;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_3;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_3;
      end
      6'b000100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_4;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_4;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_4;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_4;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_4;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_4;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_4;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_4;
      end
      6'b000101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_5;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_5;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_5;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_5;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_5;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_5;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_5;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_5;
      end
      6'b000110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_6;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_6;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_6;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_6;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_6;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_6;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_6;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_6;
      end
      6'b000111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_7;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_7;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_7;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_7;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_7;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_7;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_7;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_7;
      end
      6'b001000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_8;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_8;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_8;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_8;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_8;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_8;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_8;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_8;
      end
      6'b001001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_9;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_9;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_9;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_9;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_9;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_9;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_9;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_9;
      end
      6'b001010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_10;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_10;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_10;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_10;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_10;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_10;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_10;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_10;
      end
      6'b001011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_11;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_11;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_11;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_11;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_11;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_11;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_11;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_11;
      end
      6'b001100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_12;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_12;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_12;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_12;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_12;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_12;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_12;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_12;
      end
      6'b001101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_13;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_13;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_13;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_13;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_13;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_13;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_13;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_13;
      end
      6'b001110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_14;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_14;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_14;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_14;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_14;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_14;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_14;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_14;
      end
      6'b001111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_15;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_15;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_15;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_15;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_15;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_15;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_15;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_15;
      end
      6'b010000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_16;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_16;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_16;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_16;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_16;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_16;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_16;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_16;
      end
      6'b010001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_17;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_17;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_17;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_17;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_17;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_17;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_17;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_17;
      end
      6'b010010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_18;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_18;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_18;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_18;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_18;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_18;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_18;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_18;
      end
      6'b010011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_19;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_19;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_19;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_19;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_19;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_19;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_19;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_19;
      end
      6'b010100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_20;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_20;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_20;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_20;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_20;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_20;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_20;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_20;
      end
      6'b010101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_21;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_21;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_21;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_21;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_21;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_21;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_21;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_21;
      end
      6'b010110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_22;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_22;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_22;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_22;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_22;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_22;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_22;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_22;
      end
      6'b010111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_23;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_23;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_23;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_23;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_23;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_23;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_23;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_23;
      end
      6'b011000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_24;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_24;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_24;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_24;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_24;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_24;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_24;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_24;
      end
      6'b011001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_25;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_25;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_25;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_25;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_25;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_25;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_25;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_25;
      end
      6'b011010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_26;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_26;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_26;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_26;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_26;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_26;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_26;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_26;
      end
      6'b011011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_27;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_27;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_27;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_27;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_27;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_27;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_27;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_27;
      end
      6'b011100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_28;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_28;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_28;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_28;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_28;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_28;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_28;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_28;
      end
      6'b011101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_29;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_29;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_29;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_29;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_29;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_29;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_29;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_29;
      end
      6'b011110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_30;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_30;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_30;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_30;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_30;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_30;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_30;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_30;
      end
      6'b011111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_31;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_31;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_31;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_31;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_31;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_31;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_31;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_31;
      end
      6'b100000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_32;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_32;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_32;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_32;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_32;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_32;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_32;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_32;
      end
      6'b100001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_33;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_33;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_33;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_33;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_33;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_33;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_33;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_33;
      end
      6'b100010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_34;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_34;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_34;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_34;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_34;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_34;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_34;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_34;
      end
      6'b100011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_35;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_35;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_35;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_35;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_35;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_35;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_35;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_35;
      end
      6'b100100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_36;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_36;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_36;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_36;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_36;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_36;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_36;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_36;
      end
      6'b100101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_37;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_37;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_37;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_37;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_37;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_37;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_37;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_37;
      end
      6'b100110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_38;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_38;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_38;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_38;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_38;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_38;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_38;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_38;
      end
      6'b100111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_39;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_39;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_39;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_39;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_39;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_39;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_39;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_39;
      end
      6'b101000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_40;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_40;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_40;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_40;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_40;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_40;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_40;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_40;
      end
      6'b101001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_41;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_41;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_41;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_41;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_41;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_41;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_41;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_41;
      end
      6'b101010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_42;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_42;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_42;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_42;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_42;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_42;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_42;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_42;
      end
      6'b101011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_43;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_43;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_43;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_43;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_43;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_43;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_43;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_43;
      end
      6'b101100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_44;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_44;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_44;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_44;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_44;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_44;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_44;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_44;
      end
      6'b101101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_45;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_45;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_45;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_45;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_45;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_45;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_45;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_45;
      end
      6'b101110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_46;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_46;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_46;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_46;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_46;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_46;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_46;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_46;
      end
      6'b101111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_47;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_47;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_47;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_47;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_47;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_47;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_47;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_47;
      end
      6'b110000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_48;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_48;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_48;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_48;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_48;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_48;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_48;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_48;
      end
      6'b110001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_49;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_49;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_49;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_49;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_49;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_49;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_49;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_49;
      end
      6'b110010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_50;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_50;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_50;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_50;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_50;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_50;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_50;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_50;
      end
      6'b110011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_51;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_51;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_51;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_51;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_51;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_51;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_51;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_51;
      end
      6'b110100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_52;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_52;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_52;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_52;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_52;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_52;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_52;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_52;
      end
      6'b110101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_53;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_53;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_53;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_53;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_53;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_53;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_53;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_53;
      end
      6'b110110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_54;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_54;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_54;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_54;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_54;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_54;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_54;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_54;
      end
      6'b110111 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_55;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_55;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_55;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_55;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_55;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_55;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_55;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_55;
      end
      6'b111000 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_56;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_56;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_56;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_56;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_56;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_56;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_56;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_56;
      end
      6'b111001 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_57;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_57;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_57;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_57;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_57;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_57;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_57;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_57;
      end
      6'b111010 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_58;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_58;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_58;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_58;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_58;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_58;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_58;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_58;
      end
      6'b111011 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_59;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_59;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_59;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_59;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_59;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_59;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_59;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_59;
      end
      6'b111100 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_60;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_60;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_60;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_60;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_60;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_60;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_60;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_60;
      end
      6'b111101 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_61;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_61;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_61;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_61;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_61;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_61;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_61;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_61;
      end
      6'b111110 : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_62;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_62;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_62;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_62;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_62;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_62;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_62;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_62;
      end
      default : begin
        _zz__zz_cntRlseRespLoc_0 = cntRlseRespLoc_63;
        _zz__zz_cntLkHoldLoc_0 = cntLkHoldLoc_63;
        _zz__zz_cntLkWaitLoc_0 = cntLkWaitLoc_63;
        _zz_compLkRespLoc_getAllRlseTimeOut_1 = cntRlseRespRmt_63;
        _zz_compLkRespLoc_getAllRlseTimeOut_3 = cntLkHoldRmt_63;
        _zz_compLkRespLoc_getAllRlseTimeOut_4 = cntLkWaitRmt_63;
        _zz__zz_cntLkRespLoc_0 = cntLkRespLoc_63;
        _zz__zz_cntLkHoldWrLoc_0 = cntLkHoldWrLoc_63;
      end
    endcase
  end

  always @(*) begin
    case(compLkRespRmt_rCurTxnId)
      6'b000000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_0;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_0;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_0;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_0;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_0;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_0;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_0;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_0;
        _zz_when_TxnManCS_l261 = rAbort_0;
        _zz_when_TxnManCS_l259 = rTimeOut_0;
        _zz_when_TxnManCS_l259_1 = rReqDone_0;
      end
      6'b000001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_1;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_1;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_1;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_1;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_1;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_1;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_1;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_1;
        _zz_when_TxnManCS_l261 = rAbort_1;
        _zz_when_TxnManCS_l259 = rTimeOut_1;
        _zz_when_TxnManCS_l259_1 = rReqDone_1;
      end
      6'b000010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_2;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_2;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_2;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_2;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_2;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_2;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_2;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_2;
        _zz_when_TxnManCS_l261 = rAbort_2;
        _zz_when_TxnManCS_l259 = rTimeOut_2;
        _zz_when_TxnManCS_l259_1 = rReqDone_2;
      end
      6'b000011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_3;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_3;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_3;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_3;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_3;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_3;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_3;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_3;
        _zz_when_TxnManCS_l261 = rAbort_3;
        _zz_when_TxnManCS_l259 = rTimeOut_3;
        _zz_when_TxnManCS_l259_1 = rReqDone_3;
      end
      6'b000100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_4;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_4;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_4;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_4;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_4;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_4;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_4;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_4;
        _zz_when_TxnManCS_l261 = rAbort_4;
        _zz_when_TxnManCS_l259 = rTimeOut_4;
        _zz_when_TxnManCS_l259_1 = rReqDone_4;
      end
      6'b000101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_5;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_5;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_5;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_5;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_5;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_5;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_5;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_5;
        _zz_when_TxnManCS_l261 = rAbort_5;
        _zz_when_TxnManCS_l259 = rTimeOut_5;
        _zz_when_TxnManCS_l259_1 = rReqDone_5;
      end
      6'b000110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_6;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_6;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_6;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_6;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_6;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_6;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_6;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_6;
        _zz_when_TxnManCS_l261 = rAbort_6;
        _zz_when_TxnManCS_l259 = rTimeOut_6;
        _zz_when_TxnManCS_l259_1 = rReqDone_6;
      end
      6'b000111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_7;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_7;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_7;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_7;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_7;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_7;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_7;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_7;
        _zz_when_TxnManCS_l261 = rAbort_7;
        _zz_when_TxnManCS_l259 = rTimeOut_7;
        _zz_when_TxnManCS_l259_1 = rReqDone_7;
      end
      6'b001000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_8;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_8;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_8;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_8;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_8;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_8;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_8;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_8;
        _zz_when_TxnManCS_l261 = rAbort_8;
        _zz_when_TxnManCS_l259 = rTimeOut_8;
        _zz_when_TxnManCS_l259_1 = rReqDone_8;
      end
      6'b001001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_9;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_9;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_9;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_9;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_9;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_9;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_9;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_9;
        _zz_when_TxnManCS_l261 = rAbort_9;
        _zz_when_TxnManCS_l259 = rTimeOut_9;
        _zz_when_TxnManCS_l259_1 = rReqDone_9;
      end
      6'b001010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_10;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_10;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_10;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_10;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_10;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_10;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_10;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_10;
        _zz_when_TxnManCS_l261 = rAbort_10;
        _zz_when_TxnManCS_l259 = rTimeOut_10;
        _zz_when_TxnManCS_l259_1 = rReqDone_10;
      end
      6'b001011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_11;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_11;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_11;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_11;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_11;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_11;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_11;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_11;
        _zz_when_TxnManCS_l261 = rAbort_11;
        _zz_when_TxnManCS_l259 = rTimeOut_11;
        _zz_when_TxnManCS_l259_1 = rReqDone_11;
      end
      6'b001100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_12;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_12;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_12;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_12;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_12;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_12;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_12;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_12;
        _zz_when_TxnManCS_l261 = rAbort_12;
        _zz_when_TxnManCS_l259 = rTimeOut_12;
        _zz_when_TxnManCS_l259_1 = rReqDone_12;
      end
      6'b001101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_13;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_13;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_13;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_13;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_13;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_13;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_13;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_13;
        _zz_when_TxnManCS_l261 = rAbort_13;
        _zz_when_TxnManCS_l259 = rTimeOut_13;
        _zz_when_TxnManCS_l259_1 = rReqDone_13;
      end
      6'b001110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_14;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_14;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_14;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_14;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_14;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_14;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_14;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_14;
        _zz_when_TxnManCS_l261 = rAbort_14;
        _zz_when_TxnManCS_l259 = rTimeOut_14;
        _zz_when_TxnManCS_l259_1 = rReqDone_14;
      end
      6'b001111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_15;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_15;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_15;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_15;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_15;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_15;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_15;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_15;
        _zz_when_TxnManCS_l261 = rAbort_15;
        _zz_when_TxnManCS_l259 = rTimeOut_15;
        _zz_when_TxnManCS_l259_1 = rReqDone_15;
      end
      6'b010000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_16;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_16;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_16;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_16;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_16;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_16;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_16;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_16;
        _zz_when_TxnManCS_l261 = rAbort_16;
        _zz_when_TxnManCS_l259 = rTimeOut_16;
        _zz_when_TxnManCS_l259_1 = rReqDone_16;
      end
      6'b010001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_17;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_17;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_17;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_17;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_17;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_17;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_17;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_17;
        _zz_when_TxnManCS_l261 = rAbort_17;
        _zz_when_TxnManCS_l259 = rTimeOut_17;
        _zz_when_TxnManCS_l259_1 = rReqDone_17;
      end
      6'b010010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_18;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_18;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_18;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_18;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_18;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_18;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_18;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_18;
        _zz_when_TxnManCS_l261 = rAbort_18;
        _zz_when_TxnManCS_l259 = rTimeOut_18;
        _zz_when_TxnManCS_l259_1 = rReqDone_18;
      end
      6'b010011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_19;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_19;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_19;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_19;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_19;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_19;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_19;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_19;
        _zz_when_TxnManCS_l261 = rAbort_19;
        _zz_when_TxnManCS_l259 = rTimeOut_19;
        _zz_when_TxnManCS_l259_1 = rReqDone_19;
      end
      6'b010100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_20;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_20;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_20;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_20;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_20;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_20;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_20;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_20;
        _zz_when_TxnManCS_l261 = rAbort_20;
        _zz_when_TxnManCS_l259 = rTimeOut_20;
        _zz_when_TxnManCS_l259_1 = rReqDone_20;
      end
      6'b010101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_21;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_21;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_21;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_21;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_21;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_21;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_21;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_21;
        _zz_when_TxnManCS_l261 = rAbort_21;
        _zz_when_TxnManCS_l259 = rTimeOut_21;
        _zz_when_TxnManCS_l259_1 = rReqDone_21;
      end
      6'b010110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_22;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_22;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_22;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_22;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_22;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_22;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_22;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_22;
        _zz_when_TxnManCS_l261 = rAbort_22;
        _zz_when_TxnManCS_l259 = rTimeOut_22;
        _zz_when_TxnManCS_l259_1 = rReqDone_22;
      end
      6'b010111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_23;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_23;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_23;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_23;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_23;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_23;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_23;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_23;
        _zz_when_TxnManCS_l261 = rAbort_23;
        _zz_when_TxnManCS_l259 = rTimeOut_23;
        _zz_when_TxnManCS_l259_1 = rReqDone_23;
      end
      6'b011000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_24;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_24;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_24;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_24;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_24;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_24;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_24;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_24;
        _zz_when_TxnManCS_l261 = rAbort_24;
        _zz_when_TxnManCS_l259 = rTimeOut_24;
        _zz_when_TxnManCS_l259_1 = rReqDone_24;
      end
      6'b011001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_25;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_25;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_25;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_25;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_25;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_25;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_25;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_25;
        _zz_when_TxnManCS_l261 = rAbort_25;
        _zz_when_TxnManCS_l259 = rTimeOut_25;
        _zz_when_TxnManCS_l259_1 = rReqDone_25;
      end
      6'b011010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_26;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_26;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_26;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_26;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_26;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_26;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_26;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_26;
        _zz_when_TxnManCS_l261 = rAbort_26;
        _zz_when_TxnManCS_l259 = rTimeOut_26;
        _zz_when_TxnManCS_l259_1 = rReqDone_26;
      end
      6'b011011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_27;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_27;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_27;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_27;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_27;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_27;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_27;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_27;
        _zz_when_TxnManCS_l261 = rAbort_27;
        _zz_when_TxnManCS_l259 = rTimeOut_27;
        _zz_when_TxnManCS_l259_1 = rReqDone_27;
      end
      6'b011100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_28;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_28;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_28;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_28;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_28;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_28;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_28;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_28;
        _zz_when_TxnManCS_l261 = rAbort_28;
        _zz_when_TxnManCS_l259 = rTimeOut_28;
        _zz_when_TxnManCS_l259_1 = rReqDone_28;
      end
      6'b011101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_29;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_29;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_29;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_29;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_29;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_29;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_29;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_29;
        _zz_when_TxnManCS_l261 = rAbort_29;
        _zz_when_TxnManCS_l259 = rTimeOut_29;
        _zz_when_TxnManCS_l259_1 = rReqDone_29;
      end
      6'b011110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_30;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_30;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_30;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_30;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_30;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_30;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_30;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_30;
        _zz_when_TxnManCS_l261 = rAbort_30;
        _zz_when_TxnManCS_l259 = rTimeOut_30;
        _zz_when_TxnManCS_l259_1 = rReqDone_30;
      end
      6'b011111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_31;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_31;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_31;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_31;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_31;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_31;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_31;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_31;
        _zz_when_TxnManCS_l261 = rAbort_31;
        _zz_when_TxnManCS_l259 = rTimeOut_31;
        _zz_when_TxnManCS_l259_1 = rReqDone_31;
      end
      6'b100000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_32;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_32;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_32;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_32;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_32;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_32;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_32;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_32;
        _zz_when_TxnManCS_l261 = rAbort_32;
        _zz_when_TxnManCS_l259 = rTimeOut_32;
        _zz_when_TxnManCS_l259_1 = rReqDone_32;
      end
      6'b100001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_33;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_33;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_33;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_33;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_33;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_33;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_33;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_33;
        _zz_when_TxnManCS_l261 = rAbort_33;
        _zz_when_TxnManCS_l259 = rTimeOut_33;
        _zz_when_TxnManCS_l259_1 = rReqDone_33;
      end
      6'b100010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_34;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_34;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_34;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_34;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_34;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_34;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_34;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_34;
        _zz_when_TxnManCS_l261 = rAbort_34;
        _zz_when_TxnManCS_l259 = rTimeOut_34;
        _zz_when_TxnManCS_l259_1 = rReqDone_34;
      end
      6'b100011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_35;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_35;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_35;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_35;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_35;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_35;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_35;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_35;
        _zz_when_TxnManCS_l261 = rAbort_35;
        _zz_when_TxnManCS_l259 = rTimeOut_35;
        _zz_when_TxnManCS_l259_1 = rReqDone_35;
      end
      6'b100100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_36;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_36;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_36;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_36;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_36;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_36;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_36;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_36;
        _zz_when_TxnManCS_l261 = rAbort_36;
        _zz_when_TxnManCS_l259 = rTimeOut_36;
        _zz_when_TxnManCS_l259_1 = rReqDone_36;
      end
      6'b100101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_37;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_37;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_37;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_37;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_37;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_37;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_37;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_37;
        _zz_when_TxnManCS_l261 = rAbort_37;
        _zz_when_TxnManCS_l259 = rTimeOut_37;
        _zz_when_TxnManCS_l259_1 = rReqDone_37;
      end
      6'b100110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_38;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_38;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_38;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_38;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_38;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_38;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_38;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_38;
        _zz_when_TxnManCS_l261 = rAbort_38;
        _zz_when_TxnManCS_l259 = rTimeOut_38;
        _zz_when_TxnManCS_l259_1 = rReqDone_38;
      end
      6'b100111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_39;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_39;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_39;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_39;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_39;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_39;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_39;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_39;
        _zz_when_TxnManCS_l261 = rAbort_39;
        _zz_when_TxnManCS_l259 = rTimeOut_39;
        _zz_when_TxnManCS_l259_1 = rReqDone_39;
      end
      6'b101000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_40;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_40;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_40;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_40;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_40;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_40;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_40;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_40;
        _zz_when_TxnManCS_l261 = rAbort_40;
        _zz_when_TxnManCS_l259 = rTimeOut_40;
        _zz_when_TxnManCS_l259_1 = rReqDone_40;
      end
      6'b101001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_41;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_41;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_41;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_41;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_41;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_41;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_41;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_41;
        _zz_when_TxnManCS_l261 = rAbort_41;
        _zz_when_TxnManCS_l259 = rTimeOut_41;
        _zz_when_TxnManCS_l259_1 = rReqDone_41;
      end
      6'b101010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_42;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_42;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_42;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_42;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_42;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_42;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_42;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_42;
        _zz_when_TxnManCS_l261 = rAbort_42;
        _zz_when_TxnManCS_l259 = rTimeOut_42;
        _zz_when_TxnManCS_l259_1 = rReqDone_42;
      end
      6'b101011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_43;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_43;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_43;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_43;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_43;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_43;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_43;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_43;
        _zz_when_TxnManCS_l261 = rAbort_43;
        _zz_when_TxnManCS_l259 = rTimeOut_43;
        _zz_when_TxnManCS_l259_1 = rReqDone_43;
      end
      6'b101100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_44;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_44;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_44;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_44;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_44;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_44;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_44;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_44;
        _zz_when_TxnManCS_l261 = rAbort_44;
        _zz_when_TxnManCS_l259 = rTimeOut_44;
        _zz_when_TxnManCS_l259_1 = rReqDone_44;
      end
      6'b101101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_45;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_45;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_45;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_45;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_45;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_45;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_45;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_45;
        _zz_when_TxnManCS_l261 = rAbort_45;
        _zz_when_TxnManCS_l259 = rTimeOut_45;
        _zz_when_TxnManCS_l259_1 = rReqDone_45;
      end
      6'b101110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_46;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_46;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_46;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_46;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_46;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_46;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_46;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_46;
        _zz_when_TxnManCS_l261 = rAbort_46;
        _zz_when_TxnManCS_l259 = rTimeOut_46;
        _zz_when_TxnManCS_l259_1 = rReqDone_46;
      end
      6'b101111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_47;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_47;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_47;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_47;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_47;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_47;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_47;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_47;
        _zz_when_TxnManCS_l261 = rAbort_47;
        _zz_when_TxnManCS_l259 = rTimeOut_47;
        _zz_when_TxnManCS_l259_1 = rReqDone_47;
      end
      6'b110000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_48;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_48;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_48;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_48;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_48;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_48;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_48;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_48;
        _zz_when_TxnManCS_l261 = rAbort_48;
        _zz_when_TxnManCS_l259 = rTimeOut_48;
        _zz_when_TxnManCS_l259_1 = rReqDone_48;
      end
      6'b110001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_49;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_49;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_49;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_49;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_49;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_49;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_49;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_49;
        _zz_when_TxnManCS_l261 = rAbort_49;
        _zz_when_TxnManCS_l259 = rTimeOut_49;
        _zz_when_TxnManCS_l259_1 = rReqDone_49;
      end
      6'b110010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_50;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_50;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_50;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_50;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_50;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_50;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_50;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_50;
        _zz_when_TxnManCS_l261 = rAbort_50;
        _zz_when_TxnManCS_l259 = rTimeOut_50;
        _zz_when_TxnManCS_l259_1 = rReqDone_50;
      end
      6'b110011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_51;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_51;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_51;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_51;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_51;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_51;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_51;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_51;
        _zz_when_TxnManCS_l261 = rAbort_51;
        _zz_when_TxnManCS_l259 = rTimeOut_51;
        _zz_when_TxnManCS_l259_1 = rReqDone_51;
      end
      6'b110100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_52;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_52;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_52;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_52;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_52;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_52;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_52;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_52;
        _zz_when_TxnManCS_l261 = rAbort_52;
        _zz_when_TxnManCS_l259 = rTimeOut_52;
        _zz_when_TxnManCS_l259_1 = rReqDone_52;
      end
      6'b110101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_53;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_53;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_53;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_53;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_53;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_53;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_53;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_53;
        _zz_when_TxnManCS_l261 = rAbort_53;
        _zz_when_TxnManCS_l259 = rTimeOut_53;
        _zz_when_TxnManCS_l259_1 = rReqDone_53;
      end
      6'b110110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_54;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_54;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_54;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_54;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_54;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_54;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_54;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_54;
        _zz_when_TxnManCS_l261 = rAbort_54;
        _zz_when_TxnManCS_l259 = rTimeOut_54;
        _zz_when_TxnManCS_l259_1 = rReqDone_54;
      end
      6'b110111 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_55;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_55;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_55;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_55;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_55;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_55;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_55;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_55;
        _zz_when_TxnManCS_l261 = rAbort_55;
        _zz_when_TxnManCS_l259 = rTimeOut_55;
        _zz_when_TxnManCS_l259_1 = rReqDone_55;
      end
      6'b111000 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_56;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_56;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_56;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_56;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_56;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_56;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_56;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_56;
        _zz_when_TxnManCS_l261 = rAbort_56;
        _zz_when_TxnManCS_l259 = rTimeOut_56;
        _zz_when_TxnManCS_l259_1 = rReqDone_56;
      end
      6'b111001 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_57;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_57;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_57;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_57;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_57;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_57;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_57;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_57;
        _zz_when_TxnManCS_l261 = rAbort_57;
        _zz_when_TxnManCS_l259 = rTimeOut_57;
        _zz_when_TxnManCS_l259_1 = rReqDone_57;
      end
      6'b111010 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_58;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_58;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_58;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_58;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_58;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_58;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_58;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_58;
        _zz_when_TxnManCS_l261 = rAbort_58;
        _zz_when_TxnManCS_l259 = rTimeOut_58;
        _zz_when_TxnManCS_l259_1 = rReqDone_58;
      end
      6'b111011 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_59;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_59;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_59;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_59;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_59;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_59;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_59;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_59;
        _zz_when_TxnManCS_l261 = rAbort_59;
        _zz_when_TxnManCS_l259 = rTimeOut_59;
        _zz_when_TxnManCS_l259_1 = rReqDone_59;
      end
      6'b111100 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_60;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_60;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_60;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_60;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_60;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_60;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_60;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_60;
        _zz_when_TxnManCS_l261 = rAbort_60;
        _zz_when_TxnManCS_l259 = rTimeOut_60;
        _zz_when_TxnManCS_l259_1 = rReqDone_60;
      end
      6'b111101 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_61;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_61;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_61;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_61;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_61;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_61;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_61;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_61;
        _zz_when_TxnManCS_l261 = rAbort_61;
        _zz_when_TxnManCS_l259 = rTimeOut_61;
        _zz_when_TxnManCS_l259_1 = rReqDone_61;
      end
      6'b111110 : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_62;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_62;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_62;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_62;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_62;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_62;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_62;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_62;
        _zz_when_TxnManCS_l261 = rAbort_62;
        _zz_when_TxnManCS_l259 = rTimeOut_62;
        _zz_when_TxnManCS_l259_1 = rReqDone_62;
      end
      default : begin
        _zz_compLkRespRmt_getAllRlse = cntRlseRespLoc_63;
        _zz_compLkRespRmt_getAllRlse_1 = cntLkHoldLoc_63;
        _zz_compLkRespRmt_getAllRlse_2 = cntRlseRespRmt_63;
        _zz_compLkRespRmt_getAllRlse_3 = cntLkHoldRmt_63;
        _zz_compLkRespRmt_getAllLkResp = cntLkReqLoc_63;
        _zz_compLkRespRmt_getAllLkResp_1 = cntLkRespLoc_63;
        _zz_compLkRespRmt_getAllLkResp_2 = cntLkReqRmt_63;
        _zz_compLkRespRmt_getAllLkResp_3 = cntLkRespRmt_63;
        _zz_when_TxnManCS_l261 = rAbort_63;
        _zz_when_TxnManCS_l259 = rTimeOut_63;
        _zz_when_TxnManCS_l259_1 = rReqDone_63;
      end
    endcase
  end

  always @(*) begin
    case(io_lkRespRmt_payload_txnId)
      6'b000000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_0;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_0;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_0;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_0;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_0;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_0;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_0;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_0;
      end
      6'b000001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_1;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_1;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_1;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_1;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_1;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_1;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_1;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_1;
      end
      6'b000010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_2;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_2;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_2;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_2;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_2;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_2;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_2;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_2;
      end
      6'b000011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_3;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_3;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_3;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_3;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_3;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_3;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_3;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_3;
      end
      6'b000100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_4;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_4;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_4;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_4;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_4;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_4;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_4;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_4;
      end
      6'b000101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_5;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_5;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_5;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_5;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_5;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_5;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_5;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_5;
      end
      6'b000110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_6;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_6;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_6;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_6;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_6;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_6;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_6;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_6;
      end
      6'b000111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_7;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_7;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_7;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_7;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_7;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_7;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_7;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_7;
      end
      6'b001000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_8;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_8;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_8;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_8;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_8;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_8;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_8;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_8;
      end
      6'b001001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_9;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_9;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_9;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_9;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_9;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_9;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_9;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_9;
      end
      6'b001010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_10;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_10;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_10;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_10;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_10;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_10;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_10;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_10;
      end
      6'b001011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_11;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_11;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_11;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_11;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_11;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_11;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_11;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_11;
      end
      6'b001100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_12;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_12;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_12;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_12;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_12;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_12;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_12;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_12;
      end
      6'b001101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_13;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_13;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_13;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_13;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_13;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_13;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_13;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_13;
      end
      6'b001110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_14;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_14;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_14;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_14;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_14;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_14;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_14;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_14;
      end
      6'b001111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_15;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_15;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_15;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_15;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_15;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_15;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_15;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_15;
      end
      6'b010000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_16;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_16;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_16;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_16;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_16;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_16;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_16;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_16;
      end
      6'b010001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_17;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_17;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_17;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_17;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_17;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_17;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_17;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_17;
      end
      6'b010010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_18;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_18;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_18;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_18;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_18;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_18;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_18;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_18;
      end
      6'b010011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_19;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_19;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_19;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_19;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_19;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_19;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_19;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_19;
      end
      6'b010100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_20;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_20;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_20;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_20;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_20;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_20;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_20;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_20;
      end
      6'b010101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_21;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_21;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_21;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_21;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_21;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_21;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_21;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_21;
      end
      6'b010110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_22;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_22;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_22;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_22;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_22;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_22;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_22;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_22;
      end
      6'b010111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_23;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_23;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_23;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_23;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_23;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_23;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_23;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_23;
      end
      6'b011000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_24;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_24;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_24;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_24;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_24;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_24;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_24;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_24;
      end
      6'b011001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_25;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_25;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_25;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_25;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_25;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_25;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_25;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_25;
      end
      6'b011010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_26;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_26;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_26;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_26;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_26;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_26;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_26;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_26;
      end
      6'b011011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_27;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_27;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_27;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_27;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_27;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_27;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_27;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_27;
      end
      6'b011100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_28;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_28;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_28;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_28;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_28;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_28;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_28;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_28;
      end
      6'b011101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_29;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_29;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_29;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_29;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_29;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_29;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_29;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_29;
      end
      6'b011110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_30;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_30;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_30;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_30;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_30;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_30;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_30;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_30;
      end
      6'b011111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_31;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_31;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_31;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_31;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_31;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_31;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_31;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_31;
      end
      6'b100000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_32;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_32;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_32;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_32;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_32;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_32;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_32;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_32;
      end
      6'b100001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_33;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_33;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_33;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_33;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_33;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_33;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_33;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_33;
      end
      6'b100010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_34;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_34;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_34;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_34;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_34;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_34;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_34;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_34;
      end
      6'b100011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_35;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_35;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_35;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_35;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_35;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_35;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_35;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_35;
      end
      6'b100100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_36;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_36;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_36;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_36;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_36;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_36;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_36;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_36;
      end
      6'b100101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_37;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_37;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_37;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_37;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_37;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_37;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_37;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_37;
      end
      6'b100110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_38;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_38;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_38;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_38;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_38;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_38;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_38;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_38;
      end
      6'b100111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_39;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_39;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_39;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_39;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_39;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_39;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_39;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_39;
      end
      6'b101000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_40;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_40;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_40;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_40;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_40;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_40;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_40;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_40;
      end
      6'b101001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_41;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_41;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_41;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_41;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_41;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_41;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_41;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_41;
      end
      6'b101010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_42;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_42;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_42;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_42;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_42;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_42;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_42;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_42;
      end
      6'b101011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_43;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_43;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_43;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_43;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_43;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_43;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_43;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_43;
      end
      6'b101100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_44;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_44;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_44;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_44;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_44;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_44;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_44;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_44;
      end
      6'b101101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_45;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_45;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_45;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_45;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_45;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_45;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_45;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_45;
      end
      6'b101110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_46;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_46;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_46;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_46;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_46;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_46;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_46;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_46;
      end
      6'b101111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_47;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_47;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_47;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_47;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_47;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_47;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_47;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_47;
      end
      6'b110000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_48;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_48;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_48;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_48;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_48;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_48;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_48;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_48;
      end
      6'b110001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_49;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_49;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_49;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_49;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_49;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_49;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_49;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_49;
      end
      6'b110010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_50;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_50;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_50;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_50;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_50;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_50;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_50;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_50;
      end
      6'b110011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_51;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_51;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_51;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_51;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_51;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_51;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_51;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_51;
      end
      6'b110100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_52;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_52;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_52;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_52;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_52;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_52;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_52;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_52;
      end
      6'b110101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_53;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_53;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_53;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_53;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_53;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_53;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_53;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_53;
      end
      6'b110110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_54;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_54;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_54;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_54;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_54;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_54;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_54;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_54;
      end
      6'b110111 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_55;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_55;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_55;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_55;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_55;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_55;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_55;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_55;
      end
      6'b111000 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_56;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_56;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_56;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_56;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_56;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_56;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_56;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_56;
      end
      6'b111001 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_57;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_57;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_57;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_57;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_57;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_57;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_57;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_57;
      end
      6'b111010 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_58;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_58;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_58;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_58;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_58;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_58;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_58;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_58;
      end
      6'b111011 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_59;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_59;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_59;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_59;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_59;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_59;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_59;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_59;
      end
      6'b111100 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_60;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_60;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_60;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_60;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_60;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_60;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_60;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_60;
      end
      6'b111101 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_61;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_61;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_61;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_61;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_61;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_61;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_61;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_61;
      end
      6'b111110 : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_62;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_62;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_62;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_62;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_62;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_62;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_62;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_62;
      end
      default : begin
        _zz__zz_cntRlseRespRmt_0 = cntRlseRespRmt_63;
        _zz__zz_cntLkHoldRmt_0 = cntLkHoldRmt_63;
        _zz__zz_cntLkWaitRmt_0 = cntLkWaitRmt_63;
        _zz_compLkRespRmt_getAllRlseTimeOut = cntRlseRespLoc_63;
        _zz_compLkRespRmt_getAllRlseTimeOut_2 = cntLkHoldLoc_63;
        _zz_compLkRespRmt_getAllRlseTimeOut_3 = cntLkWaitLoc_63;
        _zz__zz_cntLkRespRmt_0 = cntLkRespRmt_63;
        _zz__zz_cntLkHoldWrRmt_0 = cntLkHoldWrRmt_63;
      end
    endcase
  end

  always @(*) begin
    case(compAxiResp_rAxiBId)
      6'b000000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_0;
      6'b000001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_1;
      6'b000010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_2;
      6'b000011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_3;
      6'b000100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_4;
      6'b000101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_5;
      6'b000110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_6;
      6'b000111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_7;
      6'b001000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_8;
      6'b001001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_9;
      6'b001010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_10;
      6'b001011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_11;
      6'b001100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_12;
      6'b001101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_13;
      6'b001110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_14;
      6'b001111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_15;
      6'b010000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_16;
      6'b010001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_17;
      6'b010010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_18;
      6'b010011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_19;
      6'b010100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_20;
      6'b010101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_21;
      6'b010110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_22;
      6'b010111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_23;
      6'b011000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_24;
      6'b011001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_25;
      6'b011010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_26;
      6'b011011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_27;
      6'b011100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_28;
      6'b011101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_29;
      6'b011110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_30;
      6'b011111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_31;
      6'b100000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_32;
      6'b100001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_33;
      6'b100010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_34;
      6'b100011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_35;
      6'b100100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_36;
      6'b100101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_37;
      6'b100110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_38;
      6'b100111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_39;
      6'b101000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_40;
      6'b101001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_41;
      6'b101010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_42;
      6'b101011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_43;
      6'b101100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_44;
      6'b101101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_45;
      6'b101110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_46;
      6'b101111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_47;
      6'b110000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_48;
      6'b110001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_49;
      6'b110010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_50;
      6'b110011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_51;
      6'b110100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_52;
      6'b110101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_53;
      6'b110110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_54;
      6'b110111 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_55;
      6'b111000 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_56;
      6'b111001 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_57;
      6'b111010 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_58;
      6'b111011 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_59;
      6'b111100 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_60;
      6'b111101 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_61;
      6'b111110 : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_62;
      default : _zz__zz_cntCmtRespLoc_0 = cntCmtRespLoc_63;
    endcase
  end

  always @(*) begin
    case(compTxnCmtLoc_curTxnId)
      6'b000000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_0;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_0;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_0;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_0;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_0;
        _zz_when_TxnManCS_l369 = rReqDone_0;
        _zz_when_TxnManCS_l369_1 = rAbort_0;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_0;
      end
      6'b000001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_1;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_1;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_1;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_1;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_1;
        _zz_when_TxnManCS_l369 = rReqDone_1;
        _zz_when_TxnManCS_l369_1 = rAbort_1;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_1;
      end
      6'b000010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_2;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_2;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_2;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_2;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_2;
        _zz_when_TxnManCS_l369 = rReqDone_2;
        _zz_when_TxnManCS_l369_1 = rAbort_2;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_2;
      end
      6'b000011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_3;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_3;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_3;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_3;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_3;
        _zz_when_TxnManCS_l369 = rReqDone_3;
        _zz_when_TxnManCS_l369_1 = rAbort_3;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_3;
      end
      6'b000100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_4;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_4;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_4;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_4;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_4;
        _zz_when_TxnManCS_l369 = rReqDone_4;
        _zz_when_TxnManCS_l369_1 = rAbort_4;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_4;
      end
      6'b000101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_5;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_5;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_5;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_5;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_5;
        _zz_when_TxnManCS_l369 = rReqDone_5;
        _zz_when_TxnManCS_l369_1 = rAbort_5;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_5;
      end
      6'b000110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_6;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_6;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_6;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_6;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_6;
        _zz_when_TxnManCS_l369 = rReqDone_6;
        _zz_when_TxnManCS_l369_1 = rAbort_6;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_6;
      end
      6'b000111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_7;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_7;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_7;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_7;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_7;
        _zz_when_TxnManCS_l369 = rReqDone_7;
        _zz_when_TxnManCS_l369_1 = rAbort_7;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_7;
      end
      6'b001000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_8;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_8;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_8;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_8;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_8;
        _zz_when_TxnManCS_l369 = rReqDone_8;
        _zz_when_TxnManCS_l369_1 = rAbort_8;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_8;
      end
      6'b001001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_9;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_9;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_9;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_9;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_9;
        _zz_when_TxnManCS_l369 = rReqDone_9;
        _zz_when_TxnManCS_l369_1 = rAbort_9;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_9;
      end
      6'b001010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_10;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_10;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_10;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_10;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_10;
        _zz_when_TxnManCS_l369 = rReqDone_10;
        _zz_when_TxnManCS_l369_1 = rAbort_10;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_10;
      end
      6'b001011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_11;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_11;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_11;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_11;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_11;
        _zz_when_TxnManCS_l369 = rReqDone_11;
        _zz_when_TxnManCS_l369_1 = rAbort_11;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_11;
      end
      6'b001100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_12;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_12;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_12;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_12;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_12;
        _zz_when_TxnManCS_l369 = rReqDone_12;
        _zz_when_TxnManCS_l369_1 = rAbort_12;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_12;
      end
      6'b001101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_13;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_13;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_13;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_13;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_13;
        _zz_when_TxnManCS_l369 = rReqDone_13;
        _zz_when_TxnManCS_l369_1 = rAbort_13;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_13;
      end
      6'b001110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_14;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_14;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_14;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_14;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_14;
        _zz_when_TxnManCS_l369 = rReqDone_14;
        _zz_when_TxnManCS_l369_1 = rAbort_14;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_14;
      end
      6'b001111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_15;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_15;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_15;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_15;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_15;
        _zz_when_TxnManCS_l369 = rReqDone_15;
        _zz_when_TxnManCS_l369_1 = rAbort_15;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_15;
      end
      6'b010000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_16;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_16;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_16;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_16;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_16;
        _zz_when_TxnManCS_l369 = rReqDone_16;
        _zz_when_TxnManCS_l369_1 = rAbort_16;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_16;
      end
      6'b010001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_17;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_17;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_17;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_17;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_17;
        _zz_when_TxnManCS_l369 = rReqDone_17;
        _zz_when_TxnManCS_l369_1 = rAbort_17;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_17;
      end
      6'b010010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_18;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_18;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_18;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_18;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_18;
        _zz_when_TxnManCS_l369 = rReqDone_18;
        _zz_when_TxnManCS_l369_1 = rAbort_18;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_18;
      end
      6'b010011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_19;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_19;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_19;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_19;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_19;
        _zz_when_TxnManCS_l369 = rReqDone_19;
        _zz_when_TxnManCS_l369_1 = rAbort_19;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_19;
      end
      6'b010100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_20;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_20;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_20;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_20;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_20;
        _zz_when_TxnManCS_l369 = rReqDone_20;
        _zz_when_TxnManCS_l369_1 = rAbort_20;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_20;
      end
      6'b010101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_21;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_21;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_21;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_21;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_21;
        _zz_when_TxnManCS_l369 = rReqDone_21;
        _zz_when_TxnManCS_l369_1 = rAbort_21;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_21;
      end
      6'b010110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_22;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_22;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_22;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_22;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_22;
        _zz_when_TxnManCS_l369 = rReqDone_22;
        _zz_when_TxnManCS_l369_1 = rAbort_22;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_22;
      end
      6'b010111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_23;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_23;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_23;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_23;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_23;
        _zz_when_TxnManCS_l369 = rReqDone_23;
        _zz_when_TxnManCS_l369_1 = rAbort_23;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_23;
      end
      6'b011000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_24;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_24;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_24;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_24;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_24;
        _zz_when_TxnManCS_l369 = rReqDone_24;
        _zz_when_TxnManCS_l369_1 = rAbort_24;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_24;
      end
      6'b011001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_25;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_25;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_25;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_25;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_25;
        _zz_when_TxnManCS_l369 = rReqDone_25;
        _zz_when_TxnManCS_l369_1 = rAbort_25;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_25;
      end
      6'b011010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_26;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_26;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_26;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_26;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_26;
        _zz_when_TxnManCS_l369 = rReqDone_26;
        _zz_when_TxnManCS_l369_1 = rAbort_26;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_26;
      end
      6'b011011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_27;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_27;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_27;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_27;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_27;
        _zz_when_TxnManCS_l369 = rReqDone_27;
        _zz_when_TxnManCS_l369_1 = rAbort_27;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_27;
      end
      6'b011100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_28;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_28;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_28;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_28;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_28;
        _zz_when_TxnManCS_l369 = rReqDone_28;
        _zz_when_TxnManCS_l369_1 = rAbort_28;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_28;
      end
      6'b011101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_29;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_29;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_29;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_29;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_29;
        _zz_when_TxnManCS_l369 = rReqDone_29;
        _zz_when_TxnManCS_l369_1 = rAbort_29;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_29;
      end
      6'b011110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_30;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_30;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_30;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_30;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_30;
        _zz_when_TxnManCS_l369 = rReqDone_30;
        _zz_when_TxnManCS_l369_1 = rAbort_30;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_30;
      end
      6'b011111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_31;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_31;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_31;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_31;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_31;
        _zz_when_TxnManCS_l369 = rReqDone_31;
        _zz_when_TxnManCS_l369_1 = rAbort_31;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_31;
      end
      6'b100000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_32;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_32;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_32;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_32;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_32;
        _zz_when_TxnManCS_l369 = rReqDone_32;
        _zz_when_TxnManCS_l369_1 = rAbort_32;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_32;
      end
      6'b100001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_33;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_33;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_33;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_33;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_33;
        _zz_when_TxnManCS_l369 = rReqDone_33;
        _zz_when_TxnManCS_l369_1 = rAbort_33;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_33;
      end
      6'b100010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_34;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_34;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_34;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_34;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_34;
        _zz_when_TxnManCS_l369 = rReqDone_34;
        _zz_when_TxnManCS_l369_1 = rAbort_34;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_34;
      end
      6'b100011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_35;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_35;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_35;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_35;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_35;
        _zz_when_TxnManCS_l369 = rReqDone_35;
        _zz_when_TxnManCS_l369_1 = rAbort_35;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_35;
      end
      6'b100100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_36;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_36;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_36;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_36;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_36;
        _zz_when_TxnManCS_l369 = rReqDone_36;
        _zz_when_TxnManCS_l369_1 = rAbort_36;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_36;
      end
      6'b100101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_37;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_37;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_37;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_37;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_37;
        _zz_when_TxnManCS_l369 = rReqDone_37;
        _zz_when_TxnManCS_l369_1 = rAbort_37;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_37;
      end
      6'b100110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_38;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_38;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_38;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_38;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_38;
        _zz_when_TxnManCS_l369 = rReqDone_38;
        _zz_when_TxnManCS_l369_1 = rAbort_38;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_38;
      end
      6'b100111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_39;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_39;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_39;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_39;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_39;
        _zz_when_TxnManCS_l369 = rReqDone_39;
        _zz_when_TxnManCS_l369_1 = rAbort_39;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_39;
      end
      6'b101000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_40;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_40;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_40;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_40;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_40;
        _zz_when_TxnManCS_l369 = rReqDone_40;
        _zz_when_TxnManCS_l369_1 = rAbort_40;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_40;
      end
      6'b101001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_41;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_41;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_41;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_41;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_41;
        _zz_when_TxnManCS_l369 = rReqDone_41;
        _zz_when_TxnManCS_l369_1 = rAbort_41;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_41;
      end
      6'b101010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_42;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_42;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_42;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_42;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_42;
        _zz_when_TxnManCS_l369 = rReqDone_42;
        _zz_when_TxnManCS_l369_1 = rAbort_42;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_42;
      end
      6'b101011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_43;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_43;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_43;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_43;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_43;
        _zz_when_TxnManCS_l369 = rReqDone_43;
        _zz_when_TxnManCS_l369_1 = rAbort_43;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_43;
      end
      6'b101100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_44;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_44;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_44;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_44;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_44;
        _zz_when_TxnManCS_l369 = rReqDone_44;
        _zz_when_TxnManCS_l369_1 = rAbort_44;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_44;
      end
      6'b101101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_45;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_45;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_45;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_45;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_45;
        _zz_when_TxnManCS_l369 = rReqDone_45;
        _zz_when_TxnManCS_l369_1 = rAbort_45;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_45;
      end
      6'b101110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_46;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_46;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_46;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_46;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_46;
        _zz_when_TxnManCS_l369 = rReqDone_46;
        _zz_when_TxnManCS_l369_1 = rAbort_46;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_46;
      end
      6'b101111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_47;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_47;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_47;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_47;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_47;
        _zz_when_TxnManCS_l369 = rReqDone_47;
        _zz_when_TxnManCS_l369_1 = rAbort_47;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_47;
      end
      6'b110000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_48;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_48;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_48;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_48;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_48;
        _zz_when_TxnManCS_l369 = rReqDone_48;
        _zz_when_TxnManCS_l369_1 = rAbort_48;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_48;
      end
      6'b110001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_49;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_49;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_49;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_49;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_49;
        _zz_when_TxnManCS_l369 = rReqDone_49;
        _zz_when_TxnManCS_l369_1 = rAbort_49;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_49;
      end
      6'b110010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_50;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_50;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_50;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_50;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_50;
        _zz_when_TxnManCS_l369 = rReqDone_50;
        _zz_when_TxnManCS_l369_1 = rAbort_50;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_50;
      end
      6'b110011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_51;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_51;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_51;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_51;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_51;
        _zz_when_TxnManCS_l369 = rReqDone_51;
        _zz_when_TxnManCS_l369_1 = rAbort_51;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_51;
      end
      6'b110100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_52;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_52;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_52;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_52;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_52;
        _zz_when_TxnManCS_l369 = rReqDone_52;
        _zz_when_TxnManCS_l369_1 = rAbort_52;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_52;
      end
      6'b110101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_53;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_53;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_53;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_53;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_53;
        _zz_when_TxnManCS_l369 = rReqDone_53;
        _zz_when_TxnManCS_l369_1 = rAbort_53;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_53;
      end
      6'b110110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_54;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_54;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_54;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_54;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_54;
        _zz_when_TxnManCS_l369 = rReqDone_54;
        _zz_when_TxnManCS_l369_1 = rAbort_54;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_54;
      end
      6'b110111 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_55;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_55;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_55;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_55;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_55;
        _zz_when_TxnManCS_l369 = rReqDone_55;
        _zz_when_TxnManCS_l369_1 = rAbort_55;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_55;
      end
      6'b111000 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_56;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_56;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_56;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_56;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_56;
        _zz_when_TxnManCS_l369 = rReqDone_56;
        _zz_when_TxnManCS_l369_1 = rAbort_56;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_56;
      end
      6'b111001 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_57;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_57;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_57;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_57;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_57;
        _zz_when_TxnManCS_l369 = rReqDone_57;
        _zz_when_TxnManCS_l369_1 = rAbort_57;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_57;
      end
      6'b111010 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_58;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_58;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_58;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_58;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_58;
        _zz_when_TxnManCS_l369 = rReqDone_58;
        _zz_when_TxnManCS_l369_1 = rAbort_58;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_58;
      end
      6'b111011 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_59;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_59;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_59;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_59;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_59;
        _zz_when_TxnManCS_l369 = rReqDone_59;
        _zz_when_TxnManCS_l369_1 = rAbort_59;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_59;
      end
      6'b111100 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_60;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_60;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_60;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_60;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_60;
        _zz_when_TxnManCS_l369 = rReqDone_60;
        _zz_when_TxnManCS_l369_1 = rAbort_60;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_60;
      end
      6'b111101 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_61;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_61;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_61;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_61;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_61;
        _zz_when_TxnManCS_l369 = rReqDone_61;
        _zz_when_TxnManCS_l369_1 = rAbort_61;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_61;
      end
      6'b111110 : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_62;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_62;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_62;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_62;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_62;
        _zz_when_TxnManCS_l369 = rReqDone_62;
        _zz_when_TxnManCS_l369_1 = rAbort_62;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_62;
      end
      default : begin
        _zz__zz_cntCmtReqLoc_0 = cntCmtReqLoc_63;
        _zz_compTxnCmtLoc_getAllLkResp = cntLkReqLoc_63;
        _zz_compTxnCmtLoc_getAllLkResp_1 = cntLkRespLoc_63;
        _zz_compTxnCmtLoc_getAllLkResp_2 = cntLkReqRmt_63;
        _zz_compTxnCmtLoc_getAllLkResp_3 = cntLkRespRmt_63;
        _zz_when_TxnManCS_l369 = rReqDone_63;
        _zz_when_TxnManCS_l369_1 = rAbort_63;
        _zz_when_TxnManCS_l369_2 = cntLkHoldWrLoc_63;
      end
    endcase
  end

  always @(*) begin
    case(compLkRlseLoc_curTxnId)
      6'b000000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_0;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_0;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_0;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_0;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_0;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_0;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_0;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_0;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_0;
        _zz_when_TxnManCS_l440_1 = rReqDone_0;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_0;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_0;
      end
      6'b000001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_1;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_1;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_1;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_1;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_1;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_1;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_1;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_1;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_1;
        _zz_when_TxnManCS_l440_1 = rReqDone_1;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_1;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_1;
      end
      6'b000010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_2;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_2;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_2;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_2;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_2;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_2;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_2;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_2;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_2;
        _zz_when_TxnManCS_l440_1 = rReqDone_2;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_2;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_2;
      end
      6'b000011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_3;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_3;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_3;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_3;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_3;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_3;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_3;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_3;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_3;
        _zz_when_TxnManCS_l440_1 = rReqDone_3;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_3;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_3;
      end
      6'b000100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_4;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_4;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_4;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_4;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_4;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_4;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_4;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_4;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_4;
        _zz_when_TxnManCS_l440_1 = rReqDone_4;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_4;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_4;
      end
      6'b000101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_5;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_5;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_5;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_5;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_5;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_5;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_5;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_5;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_5;
        _zz_when_TxnManCS_l440_1 = rReqDone_5;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_5;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_5;
      end
      6'b000110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_6;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_6;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_6;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_6;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_6;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_6;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_6;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_6;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_6;
        _zz_when_TxnManCS_l440_1 = rReqDone_6;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_6;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_6;
      end
      6'b000111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_7;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_7;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_7;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_7;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_7;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_7;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_7;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_7;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_7;
        _zz_when_TxnManCS_l440_1 = rReqDone_7;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_7;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_7;
      end
      6'b001000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_8;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_8;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_8;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_8;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_8;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_8;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_8;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_8;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_8;
        _zz_when_TxnManCS_l440_1 = rReqDone_8;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_8;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_8;
      end
      6'b001001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_9;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_9;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_9;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_9;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_9;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_9;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_9;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_9;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_9;
        _zz_when_TxnManCS_l440_1 = rReqDone_9;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_9;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_9;
      end
      6'b001010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_10;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_10;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_10;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_10;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_10;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_10;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_10;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_10;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_10;
        _zz_when_TxnManCS_l440_1 = rReqDone_10;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_10;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_10;
      end
      6'b001011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_11;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_11;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_11;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_11;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_11;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_11;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_11;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_11;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_11;
        _zz_when_TxnManCS_l440_1 = rReqDone_11;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_11;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_11;
      end
      6'b001100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_12;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_12;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_12;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_12;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_12;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_12;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_12;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_12;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_12;
        _zz_when_TxnManCS_l440_1 = rReqDone_12;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_12;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_12;
      end
      6'b001101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_13;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_13;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_13;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_13;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_13;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_13;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_13;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_13;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_13;
        _zz_when_TxnManCS_l440_1 = rReqDone_13;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_13;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_13;
      end
      6'b001110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_14;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_14;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_14;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_14;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_14;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_14;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_14;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_14;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_14;
        _zz_when_TxnManCS_l440_1 = rReqDone_14;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_14;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_14;
      end
      6'b001111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_15;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_15;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_15;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_15;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_15;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_15;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_15;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_15;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_15;
        _zz_when_TxnManCS_l440_1 = rReqDone_15;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_15;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_15;
      end
      6'b010000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_16;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_16;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_16;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_16;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_16;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_16;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_16;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_16;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_16;
        _zz_when_TxnManCS_l440_1 = rReqDone_16;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_16;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_16;
      end
      6'b010001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_17;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_17;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_17;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_17;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_17;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_17;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_17;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_17;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_17;
        _zz_when_TxnManCS_l440_1 = rReqDone_17;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_17;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_17;
      end
      6'b010010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_18;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_18;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_18;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_18;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_18;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_18;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_18;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_18;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_18;
        _zz_when_TxnManCS_l440_1 = rReqDone_18;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_18;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_18;
      end
      6'b010011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_19;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_19;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_19;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_19;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_19;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_19;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_19;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_19;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_19;
        _zz_when_TxnManCS_l440_1 = rReqDone_19;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_19;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_19;
      end
      6'b010100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_20;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_20;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_20;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_20;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_20;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_20;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_20;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_20;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_20;
        _zz_when_TxnManCS_l440_1 = rReqDone_20;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_20;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_20;
      end
      6'b010101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_21;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_21;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_21;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_21;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_21;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_21;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_21;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_21;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_21;
        _zz_when_TxnManCS_l440_1 = rReqDone_21;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_21;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_21;
      end
      6'b010110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_22;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_22;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_22;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_22;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_22;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_22;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_22;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_22;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_22;
        _zz_when_TxnManCS_l440_1 = rReqDone_22;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_22;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_22;
      end
      6'b010111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_23;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_23;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_23;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_23;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_23;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_23;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_23;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_23;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_23;
        _zz_when_TxnManCS_l440_1 = rReqDone_23;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_23;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_23;
      end
      6'b011000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_24;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_24;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_24;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_24;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_24;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_24;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_24;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_24;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_24;
        _zz_when_TxnManCS_l440_1 = rReqDone_24;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_24;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_24;
      end
      6'b011001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_25;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_25;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_25;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_25;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_25;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_25;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_25;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_25;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_25;
        _zz_when_TxnManCS_l440_1 = rReqDone_25;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_25;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_25;
      end
      6'b011010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_26;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_26;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_26;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_26;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_26;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_26;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_26;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_26;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_26;
        _zz_when_TxnManCS_l440_1 = rReqDone_26;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_26;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_26;
      end
      6'b011011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_27;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_27;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_27;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_27;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_27;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_27;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_27;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_27;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_27;
        _zz_when_TxnManCS_l440_1 = rReqDone_27;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_27;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_27;
      end
      6'b011100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_28;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_28;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_28;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_28;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_28;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_28;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_28;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_28;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_28;
        _zz_when_TxnManCS_l440_1 = rReqDone_28;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_28;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_28;
      end
      6'b011101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_29;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_29;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_29;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_29;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_29;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_29;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_29;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_29;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_29;
        _zz_when_TxnManCS_l440_1 = rReqDone_29;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_29;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_29;
      end
      6'b011110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_30;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_30;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_30;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_30;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_30;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_30;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_30;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_30;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_30;
        _zz_when_TxnManCS_l440_1 = rReqDone_30;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_30;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_30;
      end
      6'b011111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_31;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_31;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_31;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_31;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_31;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_31;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_31;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_31;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_31;
        _zz_when_TxnManCS_l440_1 = rReqDone_31;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_31;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_31;
      end
      6'b100000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_32;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_32;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_32;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_32;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_32;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_32;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_32;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_32;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_32;
        _zz_when_TxnManCS_l440_1 = rReqDone_32;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_32;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_32;
      end
      6'b100001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_33;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_33;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_33;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_33;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_33;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_33;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_33;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_33;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_33;
        _zz_when_TxnManCS_l440_1 = rReqDone_33;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_33;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_33;
      end
      6'b100010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_34;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_34;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_34;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_34;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_34;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_34;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_34;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_34;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_34;
        _zz_when_TxnManCS_l440_1 = rReqDone_34;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_34;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_34;
      end
      6'b100011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_35;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_35;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_35;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_35;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_35;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_35;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_35;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_35;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_35;
        _zz_when_TxnManCS_l440_1 = rReqDone_35;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_35;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_35;
      end
      6'b100100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_36;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_36;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_36;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_36;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_36;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_36;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_36;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_36;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_36;
        _zz_when_TxnManCS_l440_1 = rReqDone_36;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_36;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_36;
      end
      6'b100101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_37;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_37;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_37;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_37;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_37;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_37;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_37;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_37;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_37;
        _zz_when_TxnManCS_l440_1 = rReqDone_37;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_37;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_37;
      end
      6'b100110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_38;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_38;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_38;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_38;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_38;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_38;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_38;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_38;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_38;
        _zz_when_TxnManCS_l440_1 = rReqDone_38;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_38;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_38;
      end
      6'b100111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_39;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_39;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_39;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_39;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_39;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_39;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_39;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_39;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_39;
        _zz_when_TxnManCS_l440_1 = rReqDone_39;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_39;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_39;
      end
      6'b101000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_40;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_40;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_40;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_40;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_40;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_40;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_40;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_40;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_40;
        _zz_when_TxnManCS_l440_1 = rReqDone_40;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_40;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_40;
      end
      6'b101001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_41;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_41;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_41;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_41;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_41;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_41;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_41;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_41;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_41;
        _zz_when_TxnManCS_l440_1 = rReqDone_41;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_41;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_41;
      end
      6'b101010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_42;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_42;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_42;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_42;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_42;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_42;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_42;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_42;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_42;
        _zz_when_TxnManCS_l440_1 = rReqDone_42;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_42;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_42;
      end
      6'b101011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_43;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_43;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_43;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_43;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_43;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_43;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_43;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_43;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_43;
        _zz_when_TxnManCS_l440_1 = rReqDone_43;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_43;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_43;
      end
      6'b101100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_44;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_44;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_44;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_44;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_44;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_44;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_44;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_44;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_44;
        _zz_when_TxnManCS_l440_1 = rReqDone_44;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_44;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_44;
      end
      6'b101101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_45;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_45;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_45;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_45;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_45;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_45;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_45;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_45;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_45;
        _zz_when_TxnManCS_l440_1 = rReqDone_45;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_45;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_45;
      end
      6'b101110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_46;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_46;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_46;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_46;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_46;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_46;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_46;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_46;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_46;
        _zz_when_TxnManCS_l440_1 = rReqDone_46;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_46;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_46;
      end
      6'b101111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_47;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_47;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_47;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_47;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_47;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_47;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_47;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_47;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_47;
        _zz_when_TxnManCS_l440_1 = rReqDone_47;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_47;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_47;
      end
      6'b110000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_48;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_48;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_48;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_48;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_48;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_48;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_48;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_48;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_48;
        _zz_when_TxnManCS_l440_1 = rReqDone_48;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_48;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_48;
      end
      6'b110001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_49;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_49;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_49;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_49;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_49;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_49;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_49;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_49;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_49;
        _zz_when_TxnManCS_l440_1 = rReqDone_49;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_49;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_49;
      end
      6'b110010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_50;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_50;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_50;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_50;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_50;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_50;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_50;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_50;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_50;
        _zz_when_TxnManCS_l440_1 = rReqDone_50;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_50;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_50;
      end
      6'b110011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_51;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_51;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_51;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_51;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_51;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_51;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_51;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_51;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_51;
        _zz_when_TxnManCS_l440_1 = rReqDone_51;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_51;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_51;
      end
      6'b110100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_52;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_52;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_52;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_52;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_52;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_52;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_52;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_52;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_52;
        _zz_when_TxnManCS_l440_1 = rReqDone_52;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_52;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_52;
      end
      6'b110101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_53;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_53;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_53;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_53;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_53;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_53;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_53;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_53;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_53;
        _zz_when_TxnManCS_l440_1 = rReqDone_53;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_53;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_53;
      end
      6'b110110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_54;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_54;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_54;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_54;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_54;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_54;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_54;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_54;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_54;
        _zz_when_TxnManCS_l440_1 = rReqDone_54;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_54;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_54;
      end
      6'b110111 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_55;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_55;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_55;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_55;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_55;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_55;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_55;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_55;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_55;
        _zz_when_TxnManCS_l440_1 = rReqDone_55;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_55;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_55;
      end
      6'b111000 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_56;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_56;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_56;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_56;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_56;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_56;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_56;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_56;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_56;
        _zz_when_TxnManCS_l440_1 = rReqDone_56;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_56;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_56;
      end
      6'b111001 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_57;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_57;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_57;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_57;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_57;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_57;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_57;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_57;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_57;
        _zz_when_TxnManCS_l440_1 = rReqDone_57;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_57;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_57;
      end
      6'b111010 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_58;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_58;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_58;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_58;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_58;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_58;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_58;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_58;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_58;
        _zz_when_TxnManCS_l440_1 = rReqDone_58;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_58;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_58;
      end
      6'b111011 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_59;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_59;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_59;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_59;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_59;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_59;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_59;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_59;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_59;
        _zz_when_TxnManCS_l440_1 = rReqDone_59;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_59;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_59;
      end
      6'b111100 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_60;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_60;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_60;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_60;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_60;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_60;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_60;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_60;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_60;
        _zz_when_TxnManCS_l440_1 = rReqDone_60;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_60;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_60;
      end
      6'b111101 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_61;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_61;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_61;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_61;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_61;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_61;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_61;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_61;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_61;
        _zz_when_TxnManCS_l440_1 = rReqDone_61;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_61;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_61;
      end
      6'b111110 : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_62;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_62;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_62;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_62;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_62;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_62;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_62;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_62;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_62;
        _zz_when_TxnManCS_l440_1 = rReqDone_62;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_62;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_62;
      end
      default : begin
        _zz__zz_cntRlseReqLoc_0 = cntRlseReqLoc_63;
        _zz_compLkRlseLoc_getAllLkResp = cntLkReqLoc_63;
        _zz_compLkRlseLoc_getAllLkResp_1 = cntLkRespLoc_63;
        _zz_compLkRlseLoc_getAllLkResp_2 = cntLkReqRmt_63;
        _zz_compLkRlseLoc_getAllLkResp_3 = cntLkRespRmt_63;
        _zz__zz_lkReqRlseLoc_payload_txnAbt = rAbort_63;
        _zz__zz_lkReqRlseLoc_payload_txnTimeOut = rTimeOut_63;
        _zz__zz_cntRlseReqWrLoc_0 = cntRlseReqWrLoc_63;
        _zz__zz_when_TxnManCS_l440 = cntLkHoldLoc_63;
        _zz_when_TxnManCS_l440_1 = rReqDone_63;
        _zz_when_TxnManCS_l440_2 = cntCmtRespLoc_63;
        _zz_when_TxnManCS_l440_4 = cntLkWaitLoc_63;
      end
    endcase
  end

  always @(*) begin
    case(compLkRlseRmt_curTxnId)
      6'b000000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_0;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_0;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_0;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_0;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_0;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_0;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_0;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_0;
        _zz_when_TxnManCS_l489_1 = rReqDone_0;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_0;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_0;
      end
      6'b000001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_1;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_1;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_1;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_1;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_1;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_1;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_1;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_1;
        _zz_when_TxnManCS_l489_1 = rReqDone_1;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_1;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_1;
      end
      6'b000010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_2;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_2;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_2;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_2;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_2;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_2;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_2;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_2;
        _zz_when_TxnManCS_l489_1 = rReqDone_2;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_2;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_2;
      end
      6'b000011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_3;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_3;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_3;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_3;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_3;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_3;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_3;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_3;
        _zz_when_TxnManCS_l489_1 = rReqDone_3;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_3;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_3;
      end
      6'b000100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_4;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_4;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_4;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_4;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_4;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_4;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_4;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_4;
        _zz_when_TxnManCS_l489_1 = rReqDone_4;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_4;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_4;
      end
      6'b000101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_5;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_5;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_5;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_5;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_5;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_5;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_5;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_5;
        _zz_when_TxnManCS_l489_1 = rReqDone_5;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_5;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_5;
      end
      6'b000110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_6;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_6;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_6;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_6;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_6;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_6;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_6;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_6;
        _zz_when_TxnManCS_l489_1 = rReqDone_6;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_6;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_6;
      end
      6'b000111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_7;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_7;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_7;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_7;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_7;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_7;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_7;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_7;
        _zz_when_TxnManCS_l489_1 = rReqDone_7;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_7;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_7;
      end
      6'b001000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_8;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_8;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_8;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_8;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_8;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_8;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_8;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_8;
        _zz_when_TxnManCS_l489_1 = rReqDone_8;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_8;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_8;
      end
      6'b001001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_9;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_9;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_9;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_9;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_9;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_9;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_9;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_9;
        _zz_when_TxnManCS_l489_1 = rReqDone_9;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_9;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_9;
      end
      6'b001010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_10;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_10;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_10;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_10;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_10;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_10;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_10;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_10;
        _zz_when_TxnManCS_l489_1 = rReqDone_10;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_10;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_10;
      end
      6'b001011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_11;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_11;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_11;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_11;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_11;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_11;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_11;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_11;
        _zz_when_TxnManCS_l489_1 = rReqDone_11;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_11;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_11;
      end
      6'b001100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_12;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_12;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_12;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_12;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_12;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_12;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_12;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_12;
        _zz_when_TxnManCS_l489_1 = rReqDone_12;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_12;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_12;
      end
      6'b001101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_13;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_13;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_13;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_13;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_13;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_13;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_13;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_13;
        _zz_when_TxnManCS_l489_1 = rReqDone_13;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_13;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_13;
      end
      6'b001110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_14;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_14;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_14;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_14;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_14;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_14;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_14;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_14;
        _zz_when_TxnManCS_l489_1 = rReqDone_14;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_14;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_14;
      end
      6'b001111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_15;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_15;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_15;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_15;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_15;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_15;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_15;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_15;
        _zz_when_TxnManCS_l489_1 = rReqDone_15;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_15;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_15;
      end
      6'b010000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_16;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_16;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_16;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_16;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_16;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_16;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_16;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_16;
        _zz_when_TxnManCS_l489_1 = rReqDone_16;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_16;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_16;
      end
      6'b010001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_17;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_17;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_17;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_17;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_17;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_17;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_17;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_17;
        _zz_when_TxnManCS_l489_1 = rReqDone_17;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_17;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_17;
      end
      6'b010010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_18;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_18;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_18;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_18;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_18;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_18;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_18;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_18;
        _zz_when_TxnManCS_l489_1 = rReqDone_18;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_18;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_18;
      end
      6'b010011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_19;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_19;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_19;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_19;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_19;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_19;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_19;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_19;
        _zz_when_TxnManCS_l489_1 = rReqDone_19;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_19;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_19;
      end
      6'b010100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_20;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_20;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_20;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_20;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_20;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_20;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_20;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_20;
        _zz_when_TxnManCS_l489_1 = rReqDone_20;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_20;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_20;
      end
      6'b010101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_21;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_21;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_21;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_21;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_21;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_21;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_21;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_21;
        _zz_when_TxnManCS_l489_1 = rReqDone_21;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_21;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_21;
      end
      6'b010110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_22;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_22;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_22;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_22;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_22;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_22;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_22;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_22;
        _zz_when_TxnManCS_l489_1 = rReqDone_22;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_22;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_22;
      end
      6'b010111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_23;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_23;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_23;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_23;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_23;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_23;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_23;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_23;
        _zz_when_TxnManCS_l489_1 = rReqDone_23;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_23;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_23;
      end
      6'b011000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_24;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_24;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_24;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_24;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_24;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_24;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_24;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_24;
        _zz_when_TxnManCS_l489_1 = rReqDone_24;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_24;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_24;
      end
      6'b011001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_25;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_25;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_25;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_25;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_25;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_25;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_25;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_25;
        _zz_when_TxnManCS_l489_1 = rReqDone_25;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_25;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_25;
      end
      6'b011010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_26;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_26;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_26;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_26;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_26;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_26;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_26;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_26;
        _zz_when_TxnManCS_l489_1 = rReqDone_26;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_26;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_26;
      end
      6'b011011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_27;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_27;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_27;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_27;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_27;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_27;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_27;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_27;
        _zz_when_TxnManCS_l489_1 = rReqDone_27;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_27;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_27;
      end
      6'b011100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_28;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_28;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_28;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_28;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_28;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_28;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_28;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_28;
        _zz_when_TxnManCS_l489_1 = rReqDone_28;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_28;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_28;
      end
      6'b011101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_29;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_29;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_29;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_29;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_29;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_29;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_29;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_29;
        _zz_when_TxnManCS_l489_1 = rReqDone_29;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_29;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_29;
      end
      6'b011110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_30;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_30;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_30;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_30;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_30;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_30;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_30;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_30;
        _zz_when_TxnManCS_l489_1 = rReqDone_30;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_30;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_30;
      end
      6'b011111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_31;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_31;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_31;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_31;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_31;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_31;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_31;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_31;
        _zz_when_TxnManCS_l489_1 = rReqDone_31;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_31;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_31;
      end
      6'b100000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_32;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_32;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_32;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_32;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_32;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_32;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_32;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_32;
        _zz_when_TxnManCS_l489_1 = rReqDone_32;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_32;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_32;
      end
      6'b100001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_33;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_33;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_33;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_33;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_33;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_33;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_33;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_33;
        _zz_when_TxnManCS_l489_1 = rReqDone_33;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_33;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_33;
      end
      6'b100010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_34;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_34;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_34;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_34;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_34;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_34;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_34;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_34;
        _zz_when_TxnManCS_l489_1 = rReqDone_34;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_34;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_34;
      end
      6'b100011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_35;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_35;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_35;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_35;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_35;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_35;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_35;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_35;
        _zz_when_TxnManCS_l489_1 = rReqDone_35;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_35;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_35;
      end
      6'b100100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_36;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_36;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_36;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_36;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_36;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_36;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_36;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_36;
        _zz_when_TxnManCS_l489_1 = rReqDone_36;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_36;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_36;
      end
      6'b100101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_37;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_37;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_37;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_37;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_37;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_37;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_37;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_37;
        _zz_when_TxnManCS_l489_1 = rReqDone_37;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_37;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_37;
      end
      6'b100110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_38;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_38;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_38;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_38;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_38;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_38;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_38;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_38;
        _zz_when_TxnManCS_l489_1 = rReqDone_38;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_38;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_38;
      end
      6'b100111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_39;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_39;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_39;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_39;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_39;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_39;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_39;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_39;
        _zz_when_TxnManCS_l489_1 = rReqDone_39;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_39;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_39;
      end
      6'b101000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_40;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_40;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_40;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_40;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_40;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_40;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_40;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_40;
        _zz_when_TxnManCS_l489_1 = rReqDone_40;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_40;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_40;
      end
      6'b101001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_41;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_41;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_41;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_41;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_41;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_41;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_41;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_41;
        _zz_when_TxnManCS_l489_1 = rReqDone_41;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_41;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_41;
      end
      6'b101010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_42;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_42;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_42;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_42;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_42;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_42;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_42;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_42;
        _zz_when_TxnManCS_l489_1 = rReqDone_42;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_42;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_42;
      end
      6'b101011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_43;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_43;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_43;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_43;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_43;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_43;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_43;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_43;
        _zz_when_TxnManCS_l489_1 = rReqDone_43;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_43;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_43;
      end
      6'b101100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_44;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_44;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_44;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_44;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_44;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_44;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_44;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_44;
        _zz_when_TxnManCS_l489_1 = rReqDone_44;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_44;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_44;
      end
      6'b101101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_45;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_45;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_45;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_45;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_45;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_45;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_45;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_45;
        _zz_when_TxnManCS_l489_1 = rReqDone_45;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_45;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_45;
      end
      6'b101110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_46;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_46;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_46;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_46;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_46;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_46;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_46;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_46;
        _zz_when_TxnManCS_l489_1 = rReqDone_46;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_46;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_46;
      end
      6'b101111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_47;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_47;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_47;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_47;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_47;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_47;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_47;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_47;
        _zz_when_TxnManCS_l489_1 = rReqDone_47;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_47;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_47;
      end
      6'b110000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_48;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_48;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_48;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_48;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_48;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_48;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_48;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_48;
        _zz_when_TxnManCS_l489_1 = rReqDone_48;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_48;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_48;
      end
      6'b110001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_49;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_49;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_49;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_49;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_49;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_49;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_49;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_49;
        _zz_when_TxnManCS_l489_1 = rReqDone_49;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_49;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_49;
      end
      6'b110010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_50;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_50;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_50;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_50;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_50;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_50;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_50;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_50;
        _zz_when_TxnManCS_l489_1 = rReqDone_50;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_50;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_50;
      end
      6'b110011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_51;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_51;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_51;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_51;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_51;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_51;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_51;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_51;
        _zz_when_TxnManCS_l489_1 = rReqDone_51;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_51;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_51;
      end
      6'b110100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_52;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_52;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_52;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_52;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_52;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_52;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_52;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_52;
        _zz_when_TxnManCS_l489_1 = rReqDone_52;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_52;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_52;
      end
      6'b110101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_53;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_53;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_53;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_53;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_53;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_53;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_53;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_53;
        _zz_when_TxnManCS_l489_1 = rReqDone_53;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_53;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_53;
      end
      6'b110110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_54;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_54;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_54;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_54;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_54;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_54;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_54;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_54;
        _zz_when_TxnManCS_l489_1 = rReqDone_54;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_54;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_54;
      end
      6'b110111 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_55;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_55;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_55;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_55;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_55;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_55;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_55;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_55;
        _zz_when_TxnManCS_l489_1 = rReqDone_55;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_55;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_55;
      end
      6'b111000 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_56;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_56;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_56;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_56;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_56;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_56;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_56;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_56;
        _zz_when_TxnManCS_l489_1 = rReqDone_56;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_56;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_56;
      end
      6'b111001 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_57;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_57;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_57;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_57;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_57;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_57;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_57;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_57;
        _zz_when_TxnManCS_l489_1 = rReqDone_57;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_57;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_57;
      end
      6'b111010 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_58;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_58;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_58;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_58;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_58;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_58;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_58;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_58;
        _zz_when_TxnManCS_l489_1 = rReqDone_58;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_58;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_58;
      end
      6'b111011 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_59;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_59;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_59;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_59;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_59;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_59;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_59;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_59;
        _zz_when_TxnManCS_l489_1 = rReqDone_59;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_59;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_59;
      end
      6'b111100 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_60;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_60;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_60;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_60;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_60;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_60;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_60;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_60;
        _zz_when_TxnManCS_l489_1 = rReqDone_60;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_60;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_60;
      end
      6'b111101 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_61;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_61;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_61;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_61;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_61;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_61;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_61;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_61;
        _zz_when_TxnManCS_l489_1 = rReqDone_61;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_61;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_61;
      end
      6'b111110 : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_62;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_62;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_62;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_62;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_62;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_62;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_62;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_62;
        _zz_when_TxnManCS_l489_1 = rReqDone_62;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_62;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_62;
      end
      default : begin
        _zz__zz_cntRlseReqRmt_0 = cntRlseReqRmt_63;
        _zz_compLkRlseRmt_getAllLkResp = cntLkReqLoc_63;
        _zz_compLkRlseRmt_getAllLkResp_1 = cntLkRespLoc_63;
        _zz_compLkRlseRmt_getAllLkResp_2 = cntLkReqRmt_63;
        _zz_compLkRlseRmt_getAllLkResp_3 = cntLkRespRmt_63;
        _zz__zz_lkReqRlseRmt_payload_txnAbt = rAbort_63;
        _zz__zz_lkReqRlseRmt_payload_txnTimeOut = rTimeOut_63;
        _zz__zz_when_TxnManCS_l489 = cntLkHoldRmt_63;
        _zz_when_TxnManCS_l489_1 = rReqDone_63;
        _zz_when_TxnManCS_l489_3 = cntLkWaitRmt_63;
        _zz__zz_cntRlseReqWrRmt_0 = cntRlseReqWrRmt_63;
      end
    endcase
  end

  always @(*) begin
    case(compLoadTxn_cntTxnWordInLine_value)
      3'b000 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_0;
      3'b001 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_1;
      3'b010 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_2;
      3'b011 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_3;
      3'b100 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_4;
      3'b101 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_5;
      3'b110 : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_6;
      default : _zz_compLoadTxn_bitsBuff = compLoadTxn_cmdAxiDataSlice_7;
    endcase
  end

  always @(*) begin
    case(compLkReq_curTxnId)
      6'b000000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_0;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_0;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_0;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_0;
        _zz_when_TxnManCS_l128_1 = rAbort_0;
      end
      6'b000001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_1;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_1;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_1;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_1;
        _zz_when_TxnManCS_l128_1 = rAbort_1;
      end
      6'b000010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_2;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_2;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_2;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_2;
        _zz_when_TxnManCS_l128_1 = rAbort_2;
      end
      6'b000011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_3;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_3;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_3;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_3;
        _zz_when_TxnManCS_l128_1 = rAbort_3;
      end
      6'b000100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_4;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_4;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_4;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_4;
        _zz_when_TxnManCS_l128_1 = rAbort_4;
      end
      6'b000101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_5;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_5;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_5;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_5;
        _zz_when_TxnManCS_l128_1 = rAbort_5;
      end
      6'b000110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_6;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_6;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_6;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_6;
        _zz_when_TxnManCS_l128_1 = rAbort_6;
      end
      6'b000111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_7;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_7;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_7;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_7;
        _zz_when_TxnManCS_l128_1 = rAbort_7;
      end
      6'b001000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_8;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_8;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_8;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_8;
        _zz_when_TxnManCS_l128_1 = rAbort_8;
      end
      6'b001001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_9;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_9;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_9;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_9;
        _zz_when_TxnManCS_l128_1 = rAbort_9;
      end
      6'b001010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_10;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_10;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_10;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_10;
        _zz_when_TxnManCS_l128_1 = rAbort_10;
      end
      6'b001011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_11;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_11;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_11;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_11;
        _zz_when_TxnManCS_l128_1 = rAbort_11;
      end
      6'b001100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_12;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_12;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_12;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_12;
        _zz_when_TxnManCS_l128_1 = rAbort_12;
      end
      6'b001101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_13;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_13;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_13;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_13;
        _zz_when_TxnManCS_l128_1 = rAbort_13;
      end
      6'b001110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_14;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_14;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_14;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_14;
        _zz_when_TxnManCS_l128_1 = rAbort_14;
      end
      6'b001111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_15;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_15;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_15;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_15;
        _zz_when_TxnManCS_l128_1 = rAbort_15;
      end
      6'b010000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_16;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_16;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_16;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_16;
        _zz_when_TxnManCS_l128_1 = rAbort_16;
      end
      6'b010001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_17;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_17;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_17;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_17;
        _zz_when_TxnManCS_l128_1 = rAbort_17;
      end
      6'b010010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_18;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_18;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_18;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_18;
        _zz_when_TxnManCS_l128_1 = rAbort_18;
      end
      6'b010011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_19;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_19;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_19;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_19;
        _zz_when_TxnManCS_l128_1 = rAbort_19;
      end
      6'b010100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_20;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_20;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_20;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_20;
        _zz_when_TxnManCS_l128_1 = rAbort_20;
      end
      6'b010101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_21;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_21;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_21;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_21;
        _zz_when_TxnManCS_l128_1 = rAbort_21;
      end
      6'b010110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_22;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_22;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_22;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_22;
        _zz_when_TxnManCS_l128_1 = rAbort_22;
      end
      6'b010111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_23;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_23;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_23;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_23;
        _zz_when_TxnManCS_l128_1 = rAbort_23;
      end
      6'b011000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_24;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_24;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_24;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_24;
        _zz_when_TxnManCS_l128_1 = rAbort_24;
      end
      6'b011001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_25;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_25;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_25;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_25;
        _zz_when_TxnManCS_l128_1 = rAbort_25;
      end
      6'b011010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_26;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_26;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_26;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_26;
        _zz_when_TxnManCS_l128_1 = rAbort_26;
      end
      6'b011011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_27;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_27;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_27;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_27;
        _zz_when_TxnManCS_l128_1 = rAbort_27;
      end
      6'b011100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_28;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_28;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_28;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_28;
        _zz_when_TxnManCS_l128_1 = rAbort_28;
      end
      6'b011101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_29;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_29;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_29;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_29;
        _zz_when_TxnManCS_l128_1 = rAbort_29;
      end
      6'b011110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_30;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_30;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_30;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_30;
        _zz_when_TxnManCS_l128_1 = rAbort_30;
      end
      6'b011111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_31;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_31;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_31;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_31;
        _zz_when_TxnManCS_l128_1 = rAbort_31;
      end
      6'b100000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_32;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_32;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_32;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_32;
        _zz_when_TxnManCS_l128_1 = rAbort_32;
      end
      6'b100001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_33;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_33;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_33;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_33;
        _zz_when_TxnManCS_l128_1 = rAbort_33;
      end
      6'b100010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_34;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_34;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_34;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_34;
        _zz_when_TxnManCS_l128_1 = rAbort_34;
      end
      6'b100011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_35;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_35;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_35;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_35;
        _zz_when_TxnManCS_l128_1 = rAbort_35;
      end
      6'b100100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_36;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_36;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_36;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_36;
        _zz_when_TxnManCS_l128_1 = rAbort_36;
      end
      6'b100101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_37;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_37;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_37;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_37;
        _zz_when_TxnManCS_l128_1 = rAbort_37;
      end
      6'b100110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_38;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_38;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_38;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_38;
        _zz_when_TxnManCS_l128_1 = rAbort_38;
      end
      6'b100111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_39;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_39;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_39;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_39;
        _zz_when_TxnManCS_l128_1 = rAbort_39;
      end
      6'b101000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_40;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_40;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_40;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_40;
        _zz_when_TxnManCS_l128_1 = rAbort_40;
      end
      6'b101001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_41;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_41;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_41;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_41;
        _zz_when_TxnManCS_l128_1 = rAbort_41;
      end
      6'b101010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_42;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_42;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_42;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_42;
        _zz_when_TxnManCS_l128_1 = rAbort_42;
      end
      6'b101011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_43;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_43;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_43;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_43;
        _zz_when_TxnManCS_l128_1 = rAbort_43;
      end
      6'b101100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_44;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_44;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_44;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_44;
        _zz_when_TxnManCS_l128_1 = rAbort_44;
      end
      6'b101101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_45;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_45;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_45;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_45;
        _zz_when_TxnManCS_l128_1 = rAbort_45;
      end
      6'b101110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_46;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_46;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_46;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_46;
        _zz_when_TxnManCS_l128_1 = rAbort_46;
      end
      6'b101111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_47;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_47;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_47;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_47;
        _zz_when_TxnManCS_l128_1 = rAbort_47;
      end
      6'b110000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_48;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_48;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_48;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_48;
        _zz_when_TxnManCS_l128_1 = rAbort_48;
      end
      6'b110001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_49;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_49;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_49;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_49;
        _zz_when_TxnManCS_l128_1 = rAbort_49;
      end
      6'b110010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_50;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_50;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_50;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_50;
        _zz_when_TxnManCS_l128_1 = rAbort_50;
      end
      6'b110011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_51;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_51;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_51;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_51;
        _zz_when_TxnManCS_l128_1 = rAbort_51;
      end
      6'b110100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_52;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_52;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_52;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_52;
        _zz_when_TxnManCS_l128_1 = rAbort_52;
      end
      6'b110101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_53;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_53;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_53;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_53;
        _zz_when_TxnManCS_l128_1 = rAbort_53;
      end
      6'b110110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_54;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_54;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_54;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_54;
        _zz_when_TxnManCS_l128_1 = rAbort_54;
      end
      6'b110111 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_55;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_55;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_55;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_55;
        _zz_when_TxnManCS_l128_1 = rAbort_55;
      end
      6'b111000 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_56;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_56;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_56;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_56;
        _zz_when_TxnManCS_l128_1 = rAbort_56;
      end
      6'b111001 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_57;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_57;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_57;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_57;
        _zz_when_TxnManCS_l128_1 = rAbort_57;
      end
      6'b111010 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_58;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_58;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_58;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_58;
        _zz_when_TxnManCS_l128_1 = rAbort_58;
      end
      6'b111011 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_59;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_59;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_59;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_59;
        _zz_when_TxnManCS_l128_1 = rAbort_59;
      end
      6'b111100 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_60;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_60;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_60;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_60;
        _zz_when_TxnManCS_l128_1 = rAbort_60;
      end
      6'b111101 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_61;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_61;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_61;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_61;
        _zz_when_TxnManCS_l128_1 = rAbort_61;
      end
      6'b111110 : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_62;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_62;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_62;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_62;
        _zz_when_TxnManCS_l128_1 = rAbort_62;
      end
      default : begin
        _zz__zz_cntLkReqLoc_0 = cntLkReqLoc_63;
        _zz__zz_cntLkReqRmt_0 = cntLkReqRmt_63;
        _zz__zz_cntLkReqWrLoc_0 = cntLkReqWrLoc_63;
        _zz__zz_cntLkReqWrRmt_0 = cntLkReqWrRmt_63;
        _zz_when_TxnManCS_l128_1 = rAbort_63;
      end
    endcase
  end

  always @(*) begin
    case(compLoadTxn_curTxnId)
      6'b000000 : _zz_when_TxnManCS_l621 = rRlseDone_0;
      6'b000001 : _zz_when_TxnManCS_l621 = rRlseDone_1;
      6'b000010 : _zz_when_TxnManCS_l621 = rRlseDone_2;
      6'b000011 : _zz_when_TxnManCS_l621 = rRlseDone_3;
      6'b000100 : _zz_when_TxnManCS_l621 = rRlseDone_4;
      6'b000101 : _zz_when_TxnManCS_l621 = rRlseDone_5;
      6'b000110 : _zz_when_TxnManCS_l621 = rRlseDone_6;
      6'b000111 : _zz_when_TxnManCS_l621 = rRlseDone_7;
      6'b001000 : _zz_when_TxnManCS_l621 = rRlseDone_8;
      6'b001001 : _zz_when_TxnManCS_l621 = rRlseDone_9;
      6'b001010 : _zz_when_TxnManCS_l621 = rRlseDone_10;
      6'b001011 : _zz_when_TxnManCS_l621 = rRlseDone_11;
      6'b001100 : _zz_when_TxnManCS_l621 = rRlseDone_12;
      6'b001101 : _zz_when_TxnManCS_l621 = rRlseDone_13;
      6'b001110 : _zz_when_TxnManCS_l621 = rRlseDone_14;
      6'b001111 : _zz_when_TxnManCS_l621 = rRlseDone_15;
      6'b010000 : _zz_when_TxnManCS_l621 = rRlseDone_16;
      6'b010001 : _zz_when_TxnManCS_l621 = rRlseDone_17;
      6'b010010 : _zz_when_TxnManCS_l621 = rRlseDone_18;
      6'b010011 : _zz_when_TxnManCS_l621 = rRlseDone_19;
      6'b010100 : _zz_when_TxnManCS_l621 = rRlseDone_20;
      6'b010101 : _zz_when_TxnManCS_l621 = rRlseDone_21;
      6'b010110 : _zz_when_TxnManCS_l621 = rRlseDone_22;
      6'b010111 : _zz_when_TxnManCS_l621 = rRlseDone_23;
      6'b011000 : _zz_when_TxnManCS_l621 = rRlseDone_24;
      6'b011001 : _zz_when_TxnManCS_l621 = rRlseDone_25;
      6'b011010 : _zz_when_TxnManCS_l621 = rRlseDone_26;
      6'b011011 : _zz_when_TxnManCS_l621 = rRlseDone_27;
      6'b011100 : _zz_when_TxnManCS_l621 = rRlseDone_28;
      6'b011101 : _zz_when_TxnManCS_l621 = rRlseDone_29;
      6'b011110 : _zz_when_TxnManCS_l621 = rRlseDone_30;
      6'b011111 : _zz_when_TxnManCS_l621 = rRlseDone_31;
      6'b100000 : _zz_when_TxnManCS_l621 = rRlseDone_32;
      6'b100001 : _zz_when_TxnManCS_l621 = rRlseDone_33;
      6'b100010 : _zz_when_TxnManCS_l621 = rRlseDone_34;
      6'b100011 : _zz_when_TxnManCS_l621 = rRlseDone_35;
      6'b100100 : _zz_when_TxnManCS_l621 = rRlseDone_36;
      6'b100101 : _zz_when_TxnManCS_l621 = rRlseDone_37;
      6'b100110 : _zz_when_TxnManCS_l621 = rRlseDone_38;
      6'b100111 : _zz_when_TxnManCS_l621 = rRlseDone_39;
      6'b101000 : _zz_when_TxnManCS_l621 = rRlseDone_40;
      6'b101001 : _zz_when_TxnManCS_l621 = rRlseDone_41;
      6'b101010 : _zz_when_TxnManCS_l621 = rRlseDone_42;
      6'b101011 : _zz_when_TxnManCS_l621 = rRlseDone_43;
      6'b101100 : _zz_when_TxnManCS_l621 = rRlseDone_44;
      6'b101101 : _zz_when_TxnManCS_l621 = rRlseDone_45;
      6'b101110 : _zz_when_TxnManCS_l621 = rRlseDone_46;
      6'b101111 : _zz_when_TxnManCS_l621 = rRlseDone_47;
      6'b110000 : _zz_when_TxnManCS_l621 = rRlseDone_48;
      6'b110001 : _zz_when_TxnManCS_l621 = rRlseDone_49;
      6'b110010 : _zz_when_TxnManCS_l621 = rRlseDone_50;
      6'b110011 : _zz_when_TxnManCS_l621 = rRlseDone_51;
      6'b110100 : _zz_when_TxnManCS_l621 = rRlseDone_52;
      6'b110101 : _zz_when_TxnManCS_l621 = rRlseDone_53;
      6'b110110 : _zz_when_TxnManCS_l621 = rRlseDone_54;
      6'b110111 : _zz_when_TxnManCS_l621 = rRlseDone_55;
      6'b111000 : _zz_when_TxnManCS_l621 = rRlseDone_56;
      6'b111001 : _zz_when_TxnManCS_l621 = rRlseDone_57;
      6'b111010 : _zz_when_TxnManCS_l621 = rRlseDone_58;
      6'b111011 : _zz_when_TxnManCS_l621 = rRlseDone_59;
      6'b111100 : _zz_when_TxnManCS_l621 = rRlseDone_60;
      6'b111101 : _zz_when_TxnManCS_l621 = rRlseDone_61;
      6'b111110 : _zz_when_TxnManCS_l621 = rRlseDone_62;
      default : _zz_when_TxnManCS_l621 = rRlseDone_63;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReqLoc_payload_lkType)
      LkT_rd : io_lkReqLoc_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReqLoc_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReqLoc_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReqLoc_payload_lkType_string = "insTab";
      default : io_lkReqLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkReqRmt_payload_lkType)
      LkT_rd : io_lkReqRmt_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReqRmt_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReqRmt_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReqRmt_payload_lkType_string = "insTab";
      default : io_lkReqRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkRespLoc_payload_lkType)
      LkT_rd : io_lkRespLoc_payload_lkType_string = "rd    ";
      LkT_wr : io_lkRespLoc_payload_lkType_string = "wr    ";
      LkT_raw : io_lkRespLoc_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkRespLoc_payload_lkType_string = "insTab";
      default : io_lkRespLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkRespLoc_payload_respType)
      LockRespType_grant : io_lkRespLoc_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkRespLoc_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkRespLoc_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkRespLoc_payload_respType_string = "release_1";
      default : io_lkRespLoc_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_lkRespRmt_payload_lkType)
      LkT_rd : io_lkRespRmt_payload_lkType_string = "rd    ";
      LkT_wr : io_lkRespRmt_payload_lkType_string = "wr    ";
      LkT_raw : io_lkRespRmt_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkRespRmt_payload_lkType_string = "insTab";
      default : io_lkRespRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkRespRmt_payload_respType)
      LockRespType_grant : io_lkRespRmt_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkRespRmt_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkRespRmt_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkRespRmt_payload_respType_string = "release_1";
      default : io_lkRespRmt_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(lkReqGetLoc_payload_lkType)
      LkT_rd : lkReqGetLoc_payload_lkType_string = "rd    ";
      LkT_wr : lkReqGetLoc_payload_lkType_string = "wr    ";
      LkT_raw : lkReqGetLoc_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqGetLoc_payload_lkType_string = "insTab";
      default : lkReqGetLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkReqRlseLoc_payload_lkType)
      LkT_rd : lkReqRlseLoc_payload_lkType_string = "rd    ";
      LkT_wr : lkReqRlseLoc_payload_lkType_string = "wr    ";
      LkT_raw : lkReqRlseLoc_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqRlseLoc_payload_lkType_string = "insTab";
      default : lkReqRlseLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkReqGetRmt_payload_lkType)
      LkT_rd : lkReqGetRmt_payload_lkType_string = "rd    ";
      LkT_wr : lkReqGetRmt_payload_lkType_string = "wr    ";
      LkT_raw : lkReqGetRmt_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqGetRmt_payload_lkType_string = "insTab";
      default : lkReqGetRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkReqRlseRmt_payload_lkType)
      LkT_rd : lkReqRlseRmt_payload_lkType_string = "rd    ";
      LkT_wr : lkReqRlseRmt_payload_lkType_string = "wr    ";
      LkT_raw : lkReqRlseRmt_payload_lkType_string = "raw   ";
      LkT_insTab : lkReqRlseRmt_payload_lkType_string = "insTab";
      default : lkReqRlseRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_8_io_output_s2mPipe_payload_lkType)
      LkT_rd : streamArbiter_8_io_output_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamArbiter_8_io_output_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamArbiter_8_io_output_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_8_io_output_s2mPipe_payload_lkType_string = "insTab";
      default : streamArbiter_8_io_output_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_8_io_output_rData_lkType)
      LkT_rd : streamArbiter_8_io_output_rData_lkType_string = "rd    ";
      LkT_wr : streamArbiter_8_io_output_rData_lkType_string = "wr    ";
      LkT_raw : streamArbiter_8_io_output_rData_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_8_io_output_rData_lkType_string = "insTab";
      default : streamArbiter_8_io_output_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType)
      LkT_rd : _zz_payload_lkType_string = "rd    ";
      LkT_wr : _zz_payload_lkType_string = "wr    ";
      LkT_raw : _zz_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_string = "insTab";
      default : _zz_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_8_io_output_s2mPipe_rData_lkType)
      LkT_rd : streamArbiter_8_io_output_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamArbiter_8_io_output_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamArbiter_8_io_output_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_8_io_output_s2mPipe_rData_lkType_string = "insTab";
      default : streamArbiter_8_io_output_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_9_io_output_s2mPipe_payload_lkType)
      LkT_rd : streamArbiter_9_io_output_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamArbiter_9_io_output_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamArbiter_9_io_output_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_9_io_output_s2mPipe_payload_lkType_string = "insTab";
      default : streamArbiter_9_io_output_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_9_io_output_rData_lkType)
      LkT_rd : streamArbiter_9_io_output_rData_lkType_string = "rd    ";
      LkT_wr : streamArbiter_9_io_output_rData_lkType_string = "wr    ";
      LkT_raw : streamArbiter_9_io_output_rData_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_9_io_output_rData_lkType_string = "insTab";
      default : streamArbiter_9_io_output_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_1)
      LkT_rd : _zz_payload_lkType_1_string = "rd    ";
      LkT_wr : _zz_payload_lkType_1_string = "wr    ";
      LkT_raw : _zz_payload_lkType_1_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_1_string = "insTab";
      default : _zz_payload_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_9_io_output_s2mPipe_rData_lkType)
      LkT_rd : streamArbiter_9_io_output_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamArbiter_9_io_output_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamArbiter_9_io_output_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamArbiter_9_io_output_s2mPipe_rData_lkType_string = "insTab";
      default : streamArbiter_9_io_output_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkReq_txnMemRd_payload_lkType)
      LkT_rd : compLkReq_txnMemRd_payload_lkType_string = "rd    ";
      LkT_wr : compLkReq_txnMemRd_payload_lkType_string = "wr    ";
      LkT_raw : compLkReq_txnMemRd_payload_lkType_string = "raw   ";
      LkT_insTab : compLkReq_txnMemRd_payload_lkType_string = "insTab";
      default : compLkReq_txnMemRd_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkReq_txnMemRd_payload_lkType)
      LkT_rd : _zz_compLkReq_txnMemRd_payload_lkType_string = "rd    ";
      LkT_wr : _zz_compLkReq_txnMemRd_payload_lkType_string = "wr    ";
      LkT_raw : _zz_compLkReq_txnMemRd_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_compLkReq_txnMemRd_payload_lkType_string = "insTab";
      default : _zz_compLkReq_txnMemRd_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkReq_txnMemRd_payload_lkType_1)
      LkT_rd : _zz_compLkReq_txnMemRd_payload_lkType_1_string = "rd    ";
      LkT_wr : _zz_compLkReq_txnMemRd_payload_lkType_1_string = "wr    ";
      LkT_raw : _zz_compLkReq_txnMemRd_payload_lkType_1_string = "raw   ";
      LkT_insTab : _zz_compLkReq_txnMemRd_payload_lkType_1_string = "insTab";
      default : _zz_compLkReq_txnMemRd_payload_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_lkReqGetLoc_payload_lkType)
      LkT_rd : _zz_lkReqGetLoc_payload_lkType_string = "rd    ";
      LkT_wr : _zz_lkReqGetLoc_payload_lkType_string = "wr    ";
      LkT_raw : _zz_lkReqGetLoc_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_lkReqGetLoc_payload_lkType_string = "insTab";
      default : _zz_lkReqGetLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_lkReqGetRmt_payload_lkType)
      LkT_rd : _zz_lkReqGetRmt_payload_lkType_string = "rd    ";
      LkT_wr : _zz_lkReqGetRmt_payload_lkType_string = "wr    ";
      LkT_raw : _zz_lkReqGetRmt_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_lkReqGetRmt_payload_lkType_string = "insTab";
      default : _zz_lkReqGetRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRespLoc_rLkResp_payload_lkType)
      LkT_rd : compLkRespLoc_rLkResp_payload_lkType_string = "rd    ";
      LkT_wr : compLkRespLoc_rLkResp_payload_lkType_string = "wr    ";
      LkT_raw : compLkRespLoc_rLkResp_payload_lkType_string = "raw   ";
      LkT_insTab : compLkRespLoc_rLkResp_payload_lkType_string = "insTab";
      default : compLkRespLoc_rLkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRespLoc_rLkResp_payload_respType)
      LockRespType_grant : compLkRespLoc_rLkResp_payload_respType_string = "grant    ";
      LockRespType_abort : compLkRespLoc_rLkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : compLkRespLoc_rLkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : compLkRespLoc_rLkResp_payload_respType_string = "release_1";
      default : compLkRespLoc_rLkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(compLkRespRmt_rLkResp_payload_lkType)
      LkT_rd : compLkRespRmt_rLkResp_payload_lkType_string = "rd    ";
      LkT_wr : compLkRespRmt_rLkResp_payload_lkType_string = "wr    ";
      LkT_raw : compLkRespRmt_rLkResp_payload_lkType_string = "raw   ";
      LkT_insTab : compLkRespRmt_rLkResp_payload_lkType_string = "insTab";
      default : compLkRespRmt_rLkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRespRmt_rLkResp_payload_respType)
      LockRespType_grant : compLkRespRmt_rLkResp_payload_respType_string = "grant    ";
      LockRespType_abort : compLkRespRmt_rLkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : compLkRespRmt_rLkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : compLkRespRmt_rLkResp_payload_respType_string = "release_1";
      default : compLkRespRmt_rLkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(compTxnCmtLoc_cmtTxn_lkType)
      LkT_rd : compTxnCmtLoc_cmtTxn_lkType_string = "rd    ";
      LkT_wr : compTxnCmtLoc_cmtTxn_lkType_string = "wr    ";
      LkT_raw : compTxnCmtLoc_cmtTxn_lkType_string = "raw   ";
      LkT_insTab : compTxnCmtLoc_cmtTxn_lkType_string = "insTab";
      default : compTxnCmtLoc_cmtTxn_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_compTxnCmtLoc_cmtTxn_lkType)
      LkT_rd : _zz_compTxnCmtLoc_cmtTxn_lkType_string = "rd    ";
      LkT_wr : _zz_compTxnCmtLoc_cmtTxn_lkType_string = "wr    ";
      LkT_raw : _zz_compTxnCmtLoc_cmtTxn_lkType_string = "raw   ";
      LkT_insTab : _zz_compTxnCmtLoc_cmtTxn_lkType_string = "insTab";
      default : _zz_compTxnCmtLoc_cmtTxn_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compTxnCmtLoc_rCmtTxn_lkType)
      LkT_rd : compTxnCmtLoc_rCmtTxn_lkType_string = "rd    ";
      LkT_wr : compTxnCmtLoc_rCmtTxn_lkType_string = "wr    ";
      LkT_raw : compTxnCmtLoc_rCmtTxn_lkType_string = "raw   ";
      LkT_insTab : compTxnCmtLoc_rCmtTxn_lkType_string = "insTab";
      default : compTxnCmtLoc_rCmtTxn_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRlseLoc_lkItem_lkType)
      LkT_rd : compLkRlseLoc_lkItem_lkType_string = "rd    ";
      LkT_wr : compLkRlseLoc_lkItem_lkType_string = "wr    ";
      LkT_raw : compLkRlseLoc_lkItem_lkType_string = "raw   ";
      LkT_insTab : compLkRlseLoc_lkItem_lkType_string = "insTab";
      default : compLkRlseLoc_lkItem_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRlseLoc_lkItem_respType)
      LockRespType_grant : compLkRlseLoc_lkItem_respType_string = "grant    ";
      LockRespType_abort : compLkRlseLoc_lkItem_respType_string = "abort    ";
      LockRespType_waiting : compLkRlseLoc_lkItem_respType_string = "waiting  ";
      LockRespType_release_1 : compLkRlseLoc_lkItem_respType_string = "release_1";
      default : compLkRlseLoc_lkItem_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkRlseLoc_lkItem_lkType)
      LkT_rd : _zz_compLkRlseLoc_lkItem_lkType_string = "rd    ";
      LkT_wr : _zz_compLkRlseLoc_lkItem_lkType_string = "wr    ";
      LkT_raw : _zz_compLkRlseLoc_lkItem_lkType_string = "raw   ";
      LkT_insTab : _zz_compLkRlseLoc_lkItem_lkType_string = "insTab";
      default : _zz_compLkRlseLoc_lkItem_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkRlseLoc_lkItem_respType)
      LockRespType_grant : _zz_compLkRlseLoc_lkItem_respType_string = "grant    ";
      LockRespType_abort : _zz_compLkRlseLoc_lkItem_respType_string = "abort    ";
      LockRespType_waiting : _zz_compLkRlseLoc_lkItem_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_compLkRlseLoc_lkItem_respType_string = "release_1";
      default : _zz_compLkRlseLoc_lkItem_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_lkReqRlseLoc_payload_lkType)
      LkT_rd : _zz_lkReqRlseLoc_payload_lkType_string = "rd    ";
      LkT_wr : _zz_lkReqRlseLoc_payload_lkType_string = "wr    ";
      LkT_raw : _zz_lkReqRlseLoc_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_lkReqRlseLoc_payload_lkType_string = "insTab";
      default : _zz_lkReqRlseLoc_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRlseRmt_lkItem_lkType)
      LkT_rd : compLkRlseRmt_lkItem_lkType_string = "rd    ";
      LkT_wr : compLkRlseRmt_lkItem_lkType_string = "wr    ";
      LkT_raw : compLkRlseRmt_lkItem_lkType_string = "raw   ";
      LkT_insTab : compLkRlseRmt_lkItem_lkType_string = "insTab";
      default : compLkRlseRmt_lkItem_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRlseRmt_lkItem_respType)
      LockRespType_grant : compLkRlseRmt_lkItem_respType_string = "grant    ";
      LockRespType_abort : compLkRlseRmt_lkItem_respType_string = "abort    ";
      LockRespType_waiting : compLkRlseRmt_lkItem_respType_string = "waiting  ";
      LockRespType_release_1 : compLkRlseRmt_lkItem_respType_string = "release_1";
      default : compLkRlseRmt_lkItem_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkRlseRmt_lkItem_lkType)
      LkT_rd : _zz_compLkRlseRmt_lkItem_lkType_string = "rd    ";
      LkT_wr : _zz_compLkRlseRmt_lkItem_lkType_string = "wr    ";
      LkT_raw : _zz_compLkRlseRmt_lkItem_lkType_string = "raw   ";
      LkT_insTab : _zz_compLkRlseRmt_lkItem_lkType_string = "insTab";
      default : _zz_compLkRlseRmt_lkItem_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_compLkRlseRmt_lkItem_respType)
      LockRespType_grant : _zz_compLkRlseRmt_lkItem_respType_string = "grant    ";
      LockRespType_abort : _zz_compLkRlseRmt_lkItem_respType_string = "abort    ";
      LockRespType_waiting : _zz_compLkRlseRmt_lkItem_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_compLkRlseRmt_lkItem_respType_string = "release_1";
      default : _zz_compLkRlseRmt_lkItem_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_lkReqRlseRmt_payload_lkType)
      LkT_rd : _zz_lkReqRlseRmt_payload_lkType_string = "rd    ";
      LkT_wr : _zz_lkReqRlseRmt_payload_lkType_string = "wr    ";
      LkT_raw : _zz_lkReqRlseRmt_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_lkReqRlseRmt_payload_lkType_string = "insTab";
      default : _zz_lkReqRlseRmt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkReq_stateReg)
      compLkReq_enumDef_BOOT : compLkReq_stateReg_string = "BOOT  ";
      compLkReq_enumDef_CS_TXN : compLkReq_stateReg_string = "CS_TXN";
      compLkReq_enumDef_RD_TXN : compLkReq_stateReg_string = "RD_TXN";
      default : compLkReq_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkReq_stateNext)
      compLkReq_enumDef_BOOT : compLkReq_stateNext_string = "BOOT  ";
      compLkReq_enumDef_CS_TXN : compLkReq_stateNext_string = "CS_TXN";
      compLkReq_enumDef_RD_TXN : compLkReq_stateNext_string = "RD_TXN";
      default : compLkReq_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(compLkRespLoc_stateReg)
      compLkRespLoc_enumDef_BOOT : compLkRespLoc_stateReg_string = "BOOT        ";
      compLkRespLoc_enumDef_WAIT_RESP : compLkRespLoc_stateReg_string = "WAIT_RESP   ";
      compLkRespLoc_enumDef_LOCAL_RD_REQ : compLkRespLoc_stateReg_string = "LOCAL_RD_REQ";
      default : compLkRespLoc_stateReg_string = "????????????";
    endcase
  end
  always @(*) begin
    case(compLkRespLoc_stateNext)
      compLkRespLoc_enumDef_BOOT : compLkRespLoc_stateNext_string = "BOOT        ";
      compLkRespLoc_enumDef_WAIT_RESP : compLkRespLoc_stateNext_string = "WAIT_RESP   ";
      compLkRespLoc_enumDef_LOCAL_RD_REQ : compLkRespLoc_stateNext_string = "LOCAL_RD_REQ";
      default : compLkRespLoc_stateNext_string = "????????????";
    endcase
  end
  always @(*) begin
    case(compLkRespRmt_stateReg)
      compLkRespRmt_enumDef_BOOT : compLkRespRmt_stateReg_string = "BOOT          ";
      compLkRespRmt_enumDef_WAIT_RESP : compLkRespRmt_stateReg_string = "WAIT_RESP     ";
      compLkRespRmt_enumDef_RMT_RD_CONSUME : compLkRespRmt_stateReg_string = "RMT_RD_CONSUME";
      default : compLkRespRmt_stateReg_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(compLkRespRmt_stateNext)
      compLkRespRmt_enumDef_BOOT : compLkRespRmt_stateNext_string = "BOOT          ";
      compLkRespRmt_enumDef_WAIT_RESP : compLkRespRmt_stateNext_string = "WAIT_RESP     ";
      compLkRespRmt_enumDef_RMT_RD_CONSUME : compLkRespRmt_stateNext_string = "RMT_RD_CONSUME";
      default : compLkRespRmt_stateNext_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(compTxnCmtLoc_stateReg)
      compTxnCmtLoc_enumDef_BOOT : compTxnCmtLoc_stateReg_string = "BOOT    ";
      compTxnCmtLoc_enumDef_CS_TXN : compTxnCmtLoc_stateReg_string = "CS_TXN  ";
      compTxnCmtLoc_enumDef_LOCAL_AW : compTxnCmtLoc_stateReg_string = "LOCAL_AW";
      compTxnCmtLoc_enumDef_LOCAL_W : compTxnCmtLoc_stateReg_string = "LOCAL_W ";
      default : compTxnCmtLoc_stateReg_string = "????????";
    endcase
  end
  always @(*) begin
    case(compTxnCmtLoc_stateNext)
      compTxnCmtLoc_enumDef_BOOT : compTxnCmtLoc_stateNext_string = "BOOT    ";
      compTxnCmtLoc_enumDef_CS_TXN : compTxnCmtLoc_stateNext_string = "CS_TXN  ";
      compTxnCmtLoc_enumDef_LOCAL_AW : compTxnCmtLoc_stateNext_string = "LOCAL_AW";
      compTxnCmtLoc_enumDef_LOCAL_W : compTxnCmtLoc_stateNext_string = "LOCAL_W ";
      default : compTxnCmtLoc_stateNext_string = "????????";
    endcase
  end
  always @(*) begin
    case(compLkRlseLoc_stateReg)
      compLkRlseLoc_enumDef_BOOT : compLkRlseLoc_stateReg_string = "BOOT   ";
      compLkRlseLoc_enumDef_CS_TXN : compLkRlseLoc_stateReg_string = "CS_TXN ";
      compLkRlseLoc_enumDef_LK_RLSE : compLkRlseLoc_stateReg_string = "LK_RLSE";
      default : compLkRlseLoc_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(compLkRlseLoc_stateNext)
      compLkRlseLoc_enumDef_BOOT : compLkRlseLoc_stateNext_string = "BOOT   ";
      compLkRlseLoc_enumDef_CS_TXN : compLkRlseLoc_stateNext_string = "CS_TXN ";
      compLkRlseLoc_enumDef_LK_RLSE : compLkRlseLoc_stateNext_string = "LK_RLSE";
      default : compLkRlseLoc_stateNext_string = "???????";
    endcase
  end
  always @(*) begin
    case(compLkRlseRmt_stateReg)
      compLkRlseRmt_enumDef_BOOT : compLkRlseRmt_stateReg_string = "BOOT       ";
      compLkRlseRmt_enumDef_CS_TXN : compLkRlseRmt_stateReg_string = "CS_TXN     ";
      compLkRlseRmt_enumDef_RMT_LK_RLSE : compLkRlseRmt_stateReg_string = "RMT_LK_RLSE";
      compLkRlseRmt_enumDef_RMT_WR : compLkRlseRmt_stateReg_string = "RMT_WR     ";
      default : compLkRlseRmt_stateReg_string = "???????????";
    endcase
  end
  always @(*) begin
    case(compLkRlseRmt_stateNext)
      compLkRlseRmt_enumDef_BOOT : compLkRlseRmt_stateNext_string = "BOOT       ";
      compLkRlseRmt_enumDef_CS_TXN : compLkRlseRmt_stateNext_string = "CS_TXN     ";
      compLkRlseRmt_enumDef_RMT_LK_RLSE : compLkRlseRmt_stateNext_string = "RMT_LK_RLSE";
      compLkRlseRmt_enumDef_RMT_WR : compLkRlseRmt_stateNext_string = "RMT_WR     ";
      default : compLkRlseRmt_stateNext_string = "???????????";
    endcase
  end
  always @(*) begin
    case(compTimeOut_stateReg)
      compTimeOut_enumDef_BOOT : compTimeOut_stateReg_string = "BOOT ";
      compTimeOut_enumDef_IDLE : compTimeOut_stateReg_string = "IDLE ";
      compTimeOut_enumDef_COUNT : compTimeOut_stateReg_string = "COUNT";
      default : compTimeOut_stateReg_string = "?????";
    endcase
  end
  always @(*) begin
    case(compTimeOut_stateNext)
      compTimeOut_enumDef_BOOT : compTimeOut_stateNext_string = "BOOT ";
      compTimeOut_enumDef_IDLE : compTimeOut_stateNext_string = "IDLE ";
      compTimeOut_enumDef_COUNT : compTimeOut_stateNext_string = "COUNT";
      default : compTimeOut_stateNext_string = "?????";
    endcase
  end
  always @(*) begin
    case(compLoadTxn_stateReg)
      compLoadTxn_enumDef_BOOT : compLoadTxn_stateReg_string = "BOOT     ";
      compLoadTxn_enumDef_IDLE : compLoadTxn_stateReg_string = "IDLE     ";
      compLoadTxn_enumDef_CS_TXN : compLoadTxn_stateReg_string = "CS_TXN   ";
      compLoadTxn_enumDef_RD_CMDAXI : compLoadTxn_stateReg_string = "RD_CMDAXI";
      compLoadTxn_enumDef_LD_TXN : compLoadTxn_stateReg_string = "LD_TXN   ";
      default : compLoadTxn_stateReg_string = "?????????";
    endcase
  end
  always @(*) begin
    case(compLoadTxn_stateNext)
      compLoadTxn_enumDef_BOOT : compLoadTxn_stateNext_string = "BOOT     ";
      compLoadTxn_enumDef_IDLE : compLoadTxn_stateNext_string = "IDLE     ";
      compLoadTxn_enumDef_CS_TXN : compLoadTxn_stateNext_string = "CS_TXN   ";
      compLoadTxn_enumDef_RD_CMDAXI : compLoadTxn_stateNext_string = "RD_CMDAXI";
      compLoadTxn_enumDef_LD_TXN : compLoadTxn_stateNext_string = "LD_TXN   ";
      default : compLoadTxn_stateNext_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_352)
      LkT_rd : _zz_352_string = "rd    ";
      LkT_wr : _zz_352_string = "wr    ";
      LkT_raw : _zz_352_string = "raw   ";
      LkT_insTab : _zz_352_string = "insTab";
      default : _zz_352_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_353)
      LkT_rd : _zz_353_string = "rd    ";
      LkT_wr : _zz_353_string = "wr    ";
      LkT_raw : _zz_353_string = "raw   ";
      LkT_insTab : _zz_353_string = "insTab";
      default : _zz_353_string = "??????";
    endcase
  end
  always @(*) begin
    case(clkCnt_stateReg)
      clkCnt_enumDef_BOOT : clkCnt_stateReg_string = "BOOT";
      clkCnt_enumDef_IDLE : clkCnt_stateReg_string = "IDLE";
      clkCnt_enumDef_CNT : clkCnt_stateReg_string = "CNT ";
      default : clkCnt_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(clkCnt_stateNext)
      clkCnt_enumDef_BOOT : clkCnt_stateNext_string = "BOOT";
      clkCnt_enumDef_IDLE : clkCnt_stateNext_string = "IDLE";
      clkCnt_enumDef_CNT : clkCnt_stateNext_string = "CNT ";
      default : clkCnt_stateNext_string = "????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    case(compLkRespRmt_stateReg)
      compLkRespRmt_enumDef_WAIT_RESP : begin
        if(io_lkRespRmt_fire_3) begin
          if(when_TxnManCS_l303) begin
            _zz_1 = 1'b1;
          end
        end
      end
      compLkRespRmt_enumDef_RMT_RD_CONSUME : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_2 = 1'b0;
    case(compLkRespLoc_stateReg)
      compLkRespLoc_enumDef_WAIT_RESP : begin
        if(io_lkRespLoc_fire_3) begin
          if(when_TxnManCS_l214) begin
            _zz_2 = 1'b1;
          end
        end
      end
      compLkRespLoc_enumDef_LOCAL_RD_REQ : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_3 = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
      end
      compLkReq_enumDef_RD_TXN : begin
        if(compLkReq_lkReqFire) begin
          if(when_TxnManCS_l106) begin
            case(compLkReq_isLocal)
              1'b1 : begin
              end
              default : begin
                _zz_3 = 1'b1;
              end
            endcase
          end
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_4 = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
      end
      compLkReq_enumDef_RD_TXN : begin
        if(compLkReq_lkReqFire) begin
          if(when_TxnManCS_l106) begin
            case(compLkReq_isLocal)
              1'b1 : begin
                _zz_4 = 1'b1;
              end
              default : begin
              end
            endcase
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign io_cmdAxi_aw_valid = 1'b0;
  assign io_cmdAxi_w_valid = 1'b0;
  assign io_cmdAxi_aw_payload_addr = 64'h0;
  assign io_cmdAxi_aw_payload_id = 6'h0;
  assign io_cmdAxi_aw_payload_len = 8'h0;
  assign io_cmdAxi_aw_payload_size = 3'b110;
  assign io_cmdAxi_aw_payload_burst = 2'b01;
  assign io_cmdAxi_w_payload_last = 1'b0;
  assign io_cmdAxi_w_payload_data = 512'h0;
  assign io_cmdAxi_b_ready = 1'b1;
  assign io_axi_w_payload_strb = 64'hffffffffffffffff;
  assign io_cmdAxi_w_payload_strb = 64'hffffffffffffffff;
  assign lkReqGetLoc_ready = streamArbiter_8_io_inputs_0_ready;
  assign lkReqRlseLoc_ready = streamArbiter_8_io_inputs_1_ready;
  assign streamArbiter_8_io_output_ready = (! streamArbiter_8_io_output_rValid);
  assign streamArbiter_8_io_output_s2mPipe_valid = (streamArbiter_8_io_output_valid || streamArbiter_8_io_output_rValid);
  assign _zz_payload_lkType = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_lkType : streamArbiter_8_io_output_payload_lkType);
  assign streamArbiter_8_io_output_s2mPipe_payload_nId = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_nId : streamArbiter_8_io_output_payload_nId);
  assign streamArbiter_8_io_output_s2mPipe_payload_tId = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_tId : streamArbiter_8_io_output_payload_tId);
  assign streamArbiter_8_io_output_s2mPipe_payload_tabId = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_tabId : streamArbiter_8_io_output_payload_tabId);
  assign streamArbiter_8_io_output_s2mPipe_payload_snId = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_snId : streamArbiter_8_io_output_payload_snId);
  assign streamArbiter_8_io_output_s2mPipe_payload_txnId = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_txnId : streamArbiter_8_io_output_payload_txnId);
  assign streamArbiter_8_io_output_s2mPipe_payload_lkType = _zz_payload_lkType;
  assign streamArbiter_8_io_output_s2mPipe_payload_lkRelease = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_lkRelease : streamArbiter_8_io_output_payload_lkRelease);
  assign streamArbiter_8_io_output_s2mPipe_payload_txnTimeOut = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_txnTimeOut : streamArbiter_8_io_output_payload_txnTimeOut);
  assign streamArbiter_8_io_output_s2mPipe_payload_txnAbt = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_txnAbt : streamArbiter_8_io_output_payload_txnAbt);
  assign streamArbiter_8_io_output_s2mPipe_payload_lkIdx = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_lkIdx : streamArbiter_8_io_output_payload_lkIdx);
  assign streamArbiter_8_io_output_s2mPipe_payload_wLen = (streamArbiter_8_io_output_rValid ? streamArbiter_8_io_output_rData_wLen : streamArbiter_8_io_output_payload_wLen);
  always @(*) begin
    streamArbiter_8_io_output_s2mPipe_ready = streamArbiter_8_io_output_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      streamArbiter_8_io_output_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! streamArbiter_8_io_output_s2mPipe_m2sPipe_valid);
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_valid = streamArbiter_8_io_output_s2mPipe_rValid;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_nId = streamArbiter_8_io_output_s2mPipe_rData_nId;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tId = streamArbiter_8_io_output_s2mPipe_rData_tId;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tabId = streamArbiter_8_io_output_s2mPipe_rData_tabId;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_snId = streamArbiter_8_io_output_s2mPipe_rData_snId;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnId = streamArbiter_8_io_output_s2mPipe_rData_txnId;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType = streamArbiter_8_io_output_s2mPipe_rData_lkType;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkRelease = streamArbiter_8_io_output_s2mPipe_rData_lkRelease;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnTimeOut = streamArbiter_8_io_output_s2mPipe_rData_txnTimeOut;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnAbt = streamArbiter_8_io_output_s2mPipe_rData_txnAbt;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkIdx = streamArbiter_8_io_output_s2mPipe_rData_lkIdx;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_wLen = streamArbiter_8_io_output_s2mPipe_rData_wLen;
  assign io_lkReqLoc_valid = streamArbiter_8_io_output_s2mPipe_m2sPipe_valid;
  assign streamArbiter_8_io_output_s2mPipe_m2sPipe_ready = io_lkReqLoc_ready;
  assign io_lkReqLoc_payload_nId = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_nId;
  assign io_lkReqLoc_payload_tId = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tId;
  assign io_lkReqLoc_payload_tabId = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_tabId;
  assign io_lkReqLoc_payload_snId = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_snId;
  assign io_lkReqLoc_payload_txnId = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnId;
  assign io_lkReqLoc_payload_lkType = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkType;
  assign io_lkReqLoc_payload_lkRelease = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkRelease;
  assign io_lkReqLoc_payload_txnTimeOut = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnTimeOut;
  assign io_lkReqLoc_payload_txnAbt = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_txnAbt;
  assign io_lkReqLoc_payload_lkIdx = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_lkIdx;
  assign io_lkReqLoc_payload_wLen = streamArbiter_8_io_output_s2mPipe_m2sPipe_payload_wLen;
  assign lkReqGetRmt_ready = streamArbiter_9_io_inputs_0_ready;
  assign lkReqRlseRmt_ready = streamArbiter_9_io_inputs_1_ready;
  assign streamArbiter_9_io_output_ready = (! streamArbiter_9_io_output_rValid);
  assign streamArbiter_9_io_output_s2mPipe_valid = (streamArbiter_9_io_output_valid || streamArbiter_9_io_output_rValid);
  assign _zz_payload_lkType_1 = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_lkType : streamArbiter_9_io_output_payload_lkType);
  assign streamArbiter_9_io_output_s2mPipe_payload_nId = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_nId : streamArbiter_9_io_output_payload_nId);
  assign streamArbiter_9_io_output_s2mPipe_payload_tId = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_tId : streamArbiter_9_io_output_payload_tId);
  assign streamArbiter_9_io_output_s2mPipe_payload_tabId = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_tabId : streamArbiter_9_io_output_payload_tabId);
  assign streamArbiter_9_io_output_s2mPipe_payload_snId = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_snId : streamArbiter_9_io_output_payload_snId);
  assign streamArbiter_9_io_output_s2mPipe_payload_txnId = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_txnId : streamArbiter_9_io_output_payload_txnId);
  assign streamArbiter_9_io_output_s2mPipe_payload_lkType = _zz_payload_lkType_1;
  assign streamArbiter_9_io_output_s2mPipe_payload_lkRelease = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_lkRelease : streamArbiter_9_io_output_payload_lkRelease);
  assign streamArbiter_9_io_output_s2mPipe_payload_txnTimeOut = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_txnTimeOut : streamArbiter_9_io_output_payload_txnTimeOut);
  assign streamArbiter_9_io_output_s2mPipe_payload_txnAbt = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_txnAbt : streamArbiter_9_io_output_payload_txnAbt);
  assign streamArbiter_9_io_output_s2mPipe_payload_lkIdx = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_lkIdx : streamArbiter_9_io_output_payload_lkIdx);
  assign streamArbiter_9_io_output_s2mPipe_payload_wLen = (streamArbiter_9_io_output_rValid ? streamArbiter_9_io_output_rData_wLen : streamArbiter_9_io_output_payload_wLen);
  always @(*) begin
    streamArbiter_9_io_output_s2mPipe_ready = streamArbiter_9_io_output_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      streamArbiter_9_io_output_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! streamArbiter_9_io_output_s2mPipe_m2sPipe_valid);
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_valid = streamArbiter_9_io_output_s2mPipe_rValid;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_nId = streamArbiter_9_io_output_s2mPipe_rData_nId;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tId = streamArbiter_9_io_output_s2mPipe_rData_tId;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tabId = streamArbiter_9_io_output_s2mPipe_rData_tabId;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_snId = streamArbiter_9_io_output_s2mPipe_rData_snId;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnId = streamArbiter_9_io_output_s2mPipe_rData_txnId;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType = streamArbiter_9_io_output_s2mPipe_rData_lkType;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkRelease = streamArbiter_9_io_output_s2mPipe_rData_lkRelease;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnTimeOut = streamArbiter_9_io_output_s2mPipe_rData_txnTimeOut;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnAbt = streamArbiter_9_io_output_s2mPipe_rData_txnAbt;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkIdx = streamArbiter_9_io_output_s2mPipe_rData_lkIdx;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_wLen = streamArbiter_9_io_output_s2mPipe_rData_wLen;
  assign io_lkReqRmt_valid = streamArbiter_9_io_output_s2mPipe_m2sPipe_valid;
  assign streamArbiter_9_io_output_s2mPipe_m2sPipe_ready = io_lkReqRmt_ready;
  assign io_lkReqRmt_payload_nId = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_nId;
  assign io_lkReqRmt_payload_tId = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tId;
  assign io_lkReqRmt_payload_tabId = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_tabId;
  assign io_lkReqRmt_payload_snId = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_snId;
  assign io_lkReqRmt_payload_txnId = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnId;
  assign io_lkReqRmt_payload_lkType = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkType;
  assign io_lkReqRmt_payload_lkRelease = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkRelease;
  assign io_lkReqRmt_payload_txnTimeOut = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnTimeOut;
  assign io_lkReqRmt_payload_txnAbt = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_txnAbt;
  assign io_lkReqRmt_payload_lkIdx = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_lkIdx;
  assign io_lkReqRmt_payload_wLen = streamArbiter_9_io_output_s2mPipe_m2sPipe_payload_wLen;
  always @(*) begin
    lkReqGetLoc_valid = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
      end
      compLkReq_enumDef_RD_TXN : begin
        case(compLkReq_isLocal)
          1'b1 : begin
            lkReqGetLoc_valid = compLkReq_txnMemRd_valid;
          end
          default : begin
          end
        endcase
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    lkReqRlseLoc_valid = 1'b0;
    case(compLkRlseLoc_stateReg)
      compLkRlseLoc_enumDef_CS_TXN : begin
      end
      compLkRlseLoc_enumDef_LK_RLSE : begin
        lkReqRlseLoc_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    lkReqGetRmt_valid = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
      end
      compLkReq_enumDef_RD_TXN : begin
        case(compLkReq_isLocal)
          1'b1 : begin
          end
          default : begin
            lkReqGetRmt_valid = compLkReq_txnMemRd_valid;
          end
        endcase
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    lkReqRlseRmt_valid = 1'b0;
    case(compLkRlseRmt_stateReg)
      compLkRlseRmt_enumDef_CS_TXN : begin
      end
      compLkRlseRmt_enumDef_RMT_LK_RLSE : begin
        lkReqRlseRmt_valid = 1'b1;
      end
      compLkRlseRmt_enumDef_RMT_WR : begin
      end
      default : begin
      end
    endcase
  end

  assign compLkReq_wantExit = 1'b0;
  always @(*) begin
    compLkReq_wantStart = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
      end
      compLkReq_enumDef_RD_TXN : begin
      end
      default : begin
        compLkReq_wantStart = 1'b1;
      end
    endcase
  end

  assign compLkReq_wantKill = 1'b0;
  always @(*) begin
    compLkReq_txnMemRdCmd_valid = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
        if(_zz_81) begin
          compLkReq_txnMemRdCmd_valid = 1'b1;
        end
        if(compLkReq_txnMemRd_fire) begin
          compLkReq_txnMemRdCmd_valid = 1'b0;
        end
      end
      compLkReq_enumDef_RD_TXN : begin
        compLkReq_txnMemRdCmd_valid = 1'b1;
        if(when_TxnManCS_l128) begin
          compLkReq_txnMemRdCmd_valid = 1'b0;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    compLkReq_txnMemRdCmd_payload = 12'h0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
        if(_zz_81) begin
          compLkReq_txnMemRdCmd_payload = ({6'd0,compLkReq_rIdxTxn2Start} <<< 6);
        end
      end
      compLkReq_enumDef_RD_TXN : begin
        compLkReq_txnMemRdCmd_payload = (compLkReq_lkReqFire ? _zz_compLkReq_txnMemRdCmd_payload_1 : _zz_compLkReq_txnMemRdCmd_payload);
      end
      default : begin
      end
    endcase
  end

  assign _zz_compLkReq_txnMemRd_payload_nId = _zz_txnMem_port0;
  assign _zz_compLkReq_txnMemRd_payload_lkType_1 = _zz_compLkReq_txnMemRd_payload_nId[27 : 26];
  assign _zz_compLkReq_txnMemRd_payload_lkType = _zz_compLkReq_txnMemRd_payload_lkType_1;
  assign compLkReq_txnMemRd_isFree = ((! compLkReq_txnMemRd_valid) || compLkReq_txnMemRd_ready);
  assign compLkReq_txnMemRdCmd_ready = compLkReq_txnMemRd_isFree;
  assign compLkReq_txnMemRd_valid = _zz_compLkReq_txnMemRd_valid;
  assign compLkReq_txnMemRd_payload_nId = _zz_compLkReq_txnMemRd_payload_nId[0 : 0];
  assign compLkReq_txnMemRd_payload_tId = _zz_compLkReq_txnMemRd_payload_nId[22 : 1];
  assign compLkReq_txnMemRd_payload_tabId = _zz_compLkReq_txnMemRd_payload_nId[25 : 23];
  assign compLkReq_txnMemRd_payload_lkType = _zz_compLkReq_txnMemRd_payload_lkType;
  assign compLkReq_txnMemRd_payload_wLen = _zz_compLkReq_txnMemRd_payload_nId[30 : 28];
  always @(*) begin
    compLkReq_txnMemRd_ready = 1'b0;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
        if(_zz_81) begin
          compLkReq_txnMemRd_ready = 1'b1;
        end
      end
      compLkReq_enumDef_RD_TXN : begin
        compLkReq_txnMemRd_ready = compLkReq_lkReqFire;
      end
      default : begin
      end
    endcase
  end

  assign compLkReq_txnOffs = ({6'd0,compLkReq_curTxnId} <<< 6);
  assign _zz_lkReqGetLoc_payload_lkType = compLkReq_txnMemRd_payload_lkType;
  assign lkReqGetLoc_payload_nId = compLkReq_txnMemRd_payload_nId;
  assign lkReqGetLoc_payload_tId = compLkReq_txnMemRd_payload_tId;
  assign lkReqGetLoc_payload_tabId = compLkReq_txnMemRd_payload_tabId;
  assign lkReqGetLoc_payload_snId = io_nodeId;
  assign lkReqGetLoc_payload_txnId = compLkReq_curTxnId;
  assign lkReqGetLoc_payload_lkType = _zz_lkReqGetLoc_payload_lkType;
  assign lkReqGetLoc_payload_lkRelease = 1'b0;
  assign lkReqGetLoc_payload_txnTimeOut = 1'b0;
  assign lkReqGetLoc_payload_txnAbt = 1'b0;
  assign lkReqGetLoc_payload_lkIdx = compLkReq_reqIdx;
  assign lkReqGetLoc_payload_wLen = compLkReq_txnMemRd_payload_wLen;
  assign _zz_lkReqGetRmt_payload_lkType = compLkReq_txnMemRd_payload_lkType;
  assign lkReqGetRmt_payload_nId = compLkReq_txnMemRd_payload_nId;
  assign lkReqGetRmt_payload_tId = compLkReq_txnMemRd_payload_tId;
  assign lkReqGetRmt_payload_tabId = compLkReq_txnMemRd_payload_tabId;
  assign lkReqGetRmt_payload_snId = io_nodeId;
  assign lkReqGetRmt_payload_txnId = compLkReq_curTxnId;
  assign lkReqGetRmt_payload_lkType = _zz_lkReqGetRmt_payload_lkType;
  assign lkReqGetRmt_payload_lkRelease = 1'b0;
  assign lkReqGetRmt_payload_txnTimeOut = 1'b0;
  assign lkReqGetRmt_payload_txnAbt = 1'b0;
  assign lkReqGetRmt_payload_lkIdx = compLkReq_reqIdx;
  assign lkReqGetRmt_payload_wLen = compLkReq_txnMemRd_payload_wLen;
  assign compLkReq_mskTxn2Start = ((~ {rReqDone_63,{rReqDone_62,{rReqDone_61,{rReqDone_60,{_zz_compLkReq_mskTxn2Start,_zz_compLkReq_mskTxn2Start_1}}}}}) & (~ {rAbort_63,{rAbort_62,{rAbort_61,{rAbort_60,{_zz_compLkReq_mskTxn2Start_20,_zz_compLkReq_mskTxn2Start_21}}}}}));
  assign compLkReq_mskTxn2Start_ohFirst_input = compLkReq_mskTxn2Start;
  assign compLkReq_mskTxn2Start_ohFirst_masked = (compLkReq_mskTxn2Start_ohFirst_input & (~ _zz_compLkReq_mskTxn2Start_ohFirst_masked));
  assign compLkReq_mskTxn2Start_ohFirst_value = compLkReq_mskTxn2Start_ohFirst_masked;
  assign _zz_compLkReq_rIdxTxn2Start = compLkReq_mskTxn2Start_ohFirst_value[3];
  assign _zz_compLkReq_rIdxTxn2Start_1 = compLkReq_mskTxn2Start_ohFirst_value[5];
  assign _zz_compLkReq_rIdxTxn2Start_2 = compLkReq_mskTxn2Start_ohFirst_value[6];
  assign _zz_compLkReq_rIdxTxn2Start_3 = compLkReq_mskTxn2Start_ohFirst_value[7];
  assign _zz_compLkReq_rIdxTxn2Start_4 = compLkReq_mskTxn2Start_ohFirst_value[9];
  assign _zz_compLkReq_rIdxTxn2Start_5 = compLkReq_mskTxn2Start_ohFirst_value[10];
  assign _zz_compLkReq_rIdxTxn2Start_6 = compLkReq_mskTxn2Start_ohFirst_value[11];
  assign _zz_compLkReq_rIdxTxn2Start_7 = compLkReq_mskTxn2Start_ohFirst_value[12];
  assign _zz_compLkReq_rIdxTxn2Start_8 = compLkReq_mskTxn2Start_ohFirst_value[13];
  assign _zz_compLkReq_rIdxTxn2Start_9 = compLkReq_mskTxn2Start_ohFirst_value[14];
  assign _zz_compLkReq_rIdxTxn2Start_10 = compLkReq_mskTxn2Start_ohFirst_value[15];
  assign _zz_compLkReq_rIdxTxn2Start_11 = compLkReq_mskTxn2Start_ohFirst_value[17];
  assign _zz_compLkReq_rIdxTxn2Start_12 = compLkReq_mskTxn2Start_ohFirst_value[18];
  assign _zz_compLkReq_rIdxTxn2Start_13 = compLkReq_mskTxn2Start_ohFirst_value[19];
  assign _zz_compLkReq_rIdxTxn2Start_14 = compLkReq_mskTxn2Start_ohFirst_value[20];
  assign _zz_compLkReq_rIdxTxn2Start_15 = compLkReq_mskTxn2Start_ohFirst_value[21];
  assign _zz_compLkReq_rIdxTxn2Start_16 = compLkReq_mskTxn2Start_ohFirst_value[22];
  assign _zz_compLkReq_rIdxTxn2Start_17 = compLkReq_mskTxn2Start_ohFirst_value[23];
  assign _zz_compLkReq_rIdxTxn2Start_18 = compLkReq_mskTxn2Start_ohFirst_value[24];
  assign _zz_compLkReq_rIdxTxn2Start_19 = compLkReq_mskTxn2Start_ohFirst_value[25];
  assign _zz_compLkReq_rIdxTxn2Start_20 = compLkReq_mskTxn2Start_ohFirst_value[26];
  assign _zz_compLkReq_rIdxTxn2Start_21 = compLkReq_mskTxn2Start_ohFirst_value[27];
  assign _zz_compLkReq_rIdxTxn2Start_22 = compLkReq_mskTxn2Start_ohFirst_value[28];
  assign _zz_compLkReq_rIdxTxn2Start_23 = compLkReq_mskTxn2Start_ohFirst_value[29];
  assign _zz_compLkReq_rIdxTxn2Start_24 = compLkReq_mskTxn2Start_ohFirst_value[30];
  assign _zz_compLkReq_rIdxTxn2Start_25 = compLkReq_mskTxn2Start_ohFirst_value[31];
  assign _zz_compLkReq_rIdxTxn2Start_26 = compLkReq_mskTxn2Start_ohFirst_value[33];
  assign _zz_compLkReq_rIdxTxn2Start_27 = compLkReq_mskTxn2Start_ohFirst_value[34];
  assign _zz_compLkReq_rIdxTxn2Start_28 = compLkReq_mskTxn2Start_ohFirst_value[35];
  assign _zz_compLkReq_rIdxTxn2Start_29 = compLkReq_mskTxn2Start_ohFirst_value[36];
  assign _zz_compLkReq_rIdxTxn2Start_30 = compLkReq_mskTxn2Start_ohFirst_value[37];
  assign _zz_compLkReq_rIdxTxn2Start_31 = compLkReq_mskTxn2Start_ohFirst_value[38];
  assign _zz_compLkReq_rIdxTxn2Start_32 = compLkReq_mskTxn2Start_ohFirst_value[39];
  assign _zz_compLkReq_rIdxTxn2Start_33 = compLkReq_mskTxn2Start_ohFirst_value[40];
  assign _zz_compLkReq_rIdxTxn2Start_34 = compLkReq_mskTxn2Start_ohFirst_value[41];
  assign _zz_compLkReq_rIdxTxn2Start_35 = compLkReq_mskTxn2Start_ohFirst_value[42];
  assign _zz_compLkReq_rIdxTxn2Start_36 = compLkReq_mskTxn2Start_ohFirst_value[43];
  assign _zz_compLkReq_rIdxTxn2Start_37 = compLkReq_mskTxn2Start_ohFirst_value[44];
  assign _zz_compLkReq_rIdxTxn2Start_38 = compLkReq_mskTxn2Start_ohFirst_value[45];
  assign _zz_compLkReq_rIdxTxn2Start_39 = compLkReq_mskTxn2Start_ohFirst_value[46];
  assign _zz_compLkReq_rIdxTxn2Start_40 = compLkReq_mskTxn2Start_ohFirst_value[47];
  assign _zz_compLkReq_rIdxTxn2Start_41 = compLkReq_mskTxn2Start_ohFirst_value[48];
  assign _zz_compLkReq_rIdxTxn2Start_42 = compLkReq_mskTxn2Start_ohFirst_value[49];
  assign _zz_compLkReq_rIdxTxn2Start_43 = compLkReq_mskTxn2Start_ohFirst_value[50];
  assign _zz_compLkReq_rIdxTxn2Start_44 = compLkReq_mskTxn2Start_ohFirst_value[51];
  assign _zz_compLkReq_rIdxTxn2Start_45 = compLkReq_mskTxn2Start_ohFirst_value[52];
  assign _zz_compLkReq_rIdxTxn2Start_46 = compLkReq_mskTxn2Start_ohFirst_value[53];
  assign _zz_compLkReq_rIdxTxn2Start_47 = compLkReq_mskTxn2Start_ohFirst_value[54];
  assign _zz_compLkReq_rIdxTxn2Start_48 = compLkReq_mskTxn2Start_ohFirst_value[55];
  assign _zz_compLkReq_rIdxTxn2Start_49 = compLkReq_mskTxn2Start_ohFirst_value[56];
  assign _zz_compLkReq_rIdxTxn2Start_50 = compLkReq_mskTxn2Start_ohFirst_value[57];
  assign _zz_compLkReq_rIdxTxn2Start_51 = compLkReq_mskTxn2Start_ohFirst_value[58];
  assign _zz_compLkReq_rIdxTxn2Start_52 = compLkReq_mskTxn2Start_ohFirst_value[59];
  assign _zz_compLkReq_rIdxTxn2Start_53 = compLkReq_mskTxn2Start_ohFirst_value[60];
  assign _zz_compLkReq_rIdxTxn2Start_54 = compLkReq_mskTxn2Start_ohFirst_value[61];
  assign _zz_compLkReq_rIdxTxn2Start_55 = compLkReq_mskTxn2Start_ohFirst_value[62];
  assign _zz_compLkReq_rIdxTxn2Start_56 = compLkReq_mskTxn2Start_ohFirst_value[63];
  assign _zz_compLkReq_rIdxTxn2Start_57 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_57 || _zz_compLkReq_rIdxTxn2Start_26) || _zz_compLkReq_rIdxTxn2Start_28) || _zz_compLkReq_rIdxTxn2Start_30) || _zz_compLkReq_rIdxTxn2Start_32) || _zz_compLkReq_rIdxTxn2Start_34) || _zz_compLkReq_rIdxTxn2Start_36) || _zz_compLkReq_rIdxTxn2Start_38) || _zz_compLkReq_rIdxTxn2Start_40) || _zz_compLkReq_rIdxTxn2Start_42) || _zz_compLkReq_rIdxTxn2Start_44) || _zz_compLkReq_rIdxTxn2Start_46) || _zz_compLkReq_rIdxTxn2Start_48) || _zz_compLkReq_rIdxTxn2Start_50) || _zz_compLkReq_rIdxTxn2Start_52) || _zz_compLkReq_rIdxTxn2Start_54) || _zz_compLkReq_rIdxTxn2Start_56);
  assign _zz_compLkReq_rIdxTxn2Start_58 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_58 || _zz_compLkReq_rIdxTxn2Start_27) || _zz_compLkReq_rIdxTxn2Start_28) || _zz_compLkReq_rIdxTxn2Start_31) || _zz_compLkReq_rIdxTxn2Start_32) || _zz_compLkReq_rIdxTxn2Start_35) || _zz_compLkReq_rIdxTxn2Start_36) || _zz_compLkReq_rIdxTxn2Start_39) || _zz_compLkReq_rIdxTxn2Start_40) || _zz_compLkReq_rIdxTxn2Start_43) || _zz_compLkReq_rIdxTxn2Start_44) || _zz_compLkReq_rIdxTxn2Start_47) || _zz_compLkReq_rIdxTxn2Start_48) || _zz_compLkReq_rIdxTxn2Start_51) || _zz_compLkReq_rIdxTxn2Start_52) || _zz_compLkReq_rIdxTxn2Start_55) || _zz_compLkReq_rIdxTxn2Start_56);
  assign _zz_compLkReq_rIdxTxn2Start_59 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_59 || _zz_compLkReq_rIdxTxn2Start_29) || _zz_compLkReq_rIdxTxn2Start_30) || _zz_compLkReq_rIdxTxn2Start_31) || _zz_compLkReq_rIdxTxn2Start_32) || _zz_compLkReq_rIdxTxn2Start_37) || _zz_compLkReq_rIdxTxn2Start_38) || _zz_compLkReq_rIdxTxn2Start_39) || _zz_compLkReq_rIdxTxn2Start_40) || _zz_compLkReq_rIdxTxn2Start_45) || _zz_compLkReq_rIdxTxn2Start_46) || _zz_compLkReq_rIdxTxn2Start_47) || _zz_compLkReq_rIdxTxn2Start_48) || _zz_compLkReq_rIdxTxn2Start_53) || _zz_compLkReq_rIdxTxn2Start_54) || _zz_compLkReq_rIdxTxn2Start_55) || _zz_compLkReq_rIdxTxn2Start_56);
  assign _zz_compLkReq_rIdxTxn2Start_60 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_60 || _zz_compLkReq_rIdxTxn2Start_33) || _zz_compLkReq_rIdxTxn2Start_34) || _zz_compLkReq_rIdxTxn2Start_35) || _zz_compLkReq_rIdxTxn2Start_36) || _zz_compLkReq_rIdxTxn2Start_37) || _zz_compLkReq_rIdxTxn2Start_38) || _zz_compLkReq_rIdxTxn2Start_39) || _zz_compLkReq_rIdxTxn2Start_40) || _zz_compLkReq_rIdxTxn2Start_49) || _zz_compLkReq_rIdxTxn2Start_50) || _zz_compLkReq_rIdxTxn2Start_51) || _zz_compLkReq_rIdxTxn2Start_52) || _zz_compLkReq_rIdxTxn2Start_53) || _zz_compLkReq_rIdxTxn2Start_54) || _zz_compLkReq_rIdxTxn2Start_55) || _zz_compLkReq_rIdxTxn2Start_56);
  assign _zz_compLkReq_rIdxTxn2Start_61 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_61 || _zz_compLkReq_rIdxTxn2Start_41) || _zz_compLkReq_rIdxTxn2Start_42) || _zz_compLkReq_rIdxTxn2Start_43) || _zz_compLkReq_rIdxTxn2Start_44) || _zz_compLkReq_rIdxTxn2Start_45) || _zz_compLkReq_rIdxTxn2Start_46) || _zz_compLkReq_rIdxTxn2Start_47) || _zz_compLkReq_rIdxTxn2Start_48) || _zz_compLkReq_rIdxTxn2Start_49) || _zz_compLkReq_rIdxTxn2Start_50) || _zz_compLkReq_rIdxTxn2Start_51) || _zz_compLkReq_rIdxTxn2Start_52) || _zz_compLkReq_rIdxTxn2Start_53) || _zz_compLkReq_rIdxTxn2Start_54) || _zz_compLkReq_rIdxTxn2Start_55) || _zz_compLkReq_rIdxTxn2Start_56);
  assign _zz_compLkReq_rIdxTxn2Start_62 = ((((((((((((((((_zz__zz_compLkReq_rIdxTxn2Start_62 || _zz_compLkReq_rIdxTxn2Start_41) || _zz_compLkReq_rIdxTxn2Start_42) || _zz_compLkReq_rIdxTxn2Start_43) || _zz_compLkReq_rIdxTxn2Start_44) || _zz_compLkReq_rIdxTxn2Start_45) || _zz_compLkReq_rIdxTxn2Start_46) || _zz_compLkReq_rIdxTxn2Start_47) || _zz_compLkReq_rIdxTxn2Start_48) || _zz_compLkReq_rIdxTxn2Start_49) || _zz_compLkReq_rIdxTxn2Start_50) || _zz_compLkReq_rIdxTxn2Start_51) || _zz_compLkReq_rIdxTxn2Start_52) || _zz_compLkReq_rIdxTxn2Start_53) || _zz_compLkReq_rIdxTxn2Start_54) || _zz_compLkReq_rIdxTxn2Start_55) || _zz_compLkReq_rIdxTxn2Start_56);
  assign lkReqGetLoc_fire = (lkReqGetLoc_valid && lkReqGetLoc_ready);
  assign lkReqGetRmt_fire = (lkReqGetRmt_valid && lkReqGetRmt_ready);
  assign compLkReq_lkReqFire = (lkReqGetLoc_fire || lkReqGetRmt_fire);
  assign compLkReq_isLocal = (compLkReq_txnMemRd_payload_nId == io_nodeId);
  assign compLkRespLoc_wantExit = 1'b0;
  always @(*) begin
    compLkRespLoc_wantStart = 1'b0;
    case(compLkRespLoc_stateReg)
      compLkRespLoc_enumDef_WAIT_RESP : begin
      end
      compLkRespLoc_enumDef_LOCAL_RD_REQ : begin
      end
      default : begin
        compLkRespLoc_wantStart = 1'b1;
      end
    endcase
  end

  assign compLkRespLoc_wantKill = 1'b0;
  assign io_lkRespLoc_fire = (io_lkRespLoc_valid && io_lkRespLoc_ready);
  assign compLkRespLoc_txnOffs = ({6'd0,io_lkRespLoc_payload_txnId} <<< 6);
  assign io_lkRespLoc_fire_1 = (io_lkRespLoc_valid && io_lkRespLoc_ready);
  assign compLkRespLoc_getAllRlse = ((_zz_compLkRespLoc_getAllRlse == _zz_compLkRespLoc_getAllRlse_1) && (_zz_compLkRespLoc_getAllRlse_2 == _zz_compLkRespLoc_getAllRlse_3));
  assign compLkRespLoc_getAllLkResp = ((_zz_compLkRespLoc_getAllLkResp == _zz_compLkRespLoc_getAllLkResp_1) && (_zz_compLkRespLoc_getAllLkResp_2 == _zz_compLkRespLoc_getAllLkResp_3));
  assign _zz_cntRlseRespLoc_0 = _zz__zz_cntRlseRespLoc_0;
  assign _zz_5 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign _zz_cntLkHoldLoc_0 = _zz__zz_cntLkHoldLoc_0;
  assign _zz_6 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign _zz_cntLkWaitLoc_0 = _zz__zz_cntLkWaitLoc_0;
  assign _zz_7 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign compLkRespLoc_getAllRlseTimeOut = ((_zz_cntRlseRespLoc_0 == _zz_compLkRespLoc_getAllRlseTimeOut) && (_zz_compLkRespLoc_getAllRlseTimeOut_1 == _zz_compLkRespLoc_getAllRlseTimeOut_2));
  assign when_TxnManCS_l166 = _zz_when_TxnManCS_l166;
  assign io_lkReqLoc_fire = (io_lkReqLoc_valid && io_lkReqLoc_ready);
  assign io_lkReqRmt_fire = (io_lkReqRmt_valid && io_lkReqRmt_ready);
  assign compLkRespLoc_firstReqAbt = ((when_TxnManCS_l166 && (! (io_lkReqLoc_fire && (io_lkReqLoc_payload_txnId == compLkRespLoc_rCurTxnId)))) && (! (io_lkReqRmt_fire && (io_lkReqRmt_payload_txnId == compLkRespLoc_rCurTxnId))));
  assign io_lkRespLoc_fire_2 = (io_lkRespLoc_valid && io_lkRespLoc_ready);
  assign when_TxnManCS_l164 = ((compLkRespLoc_rFire && ((compLkRespLoc_getAllRlse && compLkRespLoc_getAllLkResp) || (_zz_when_TxnManCS_l164 && compLkRespLoc_getAllRlseTimeOut))) && (_zz_when_TxnManCS_l164_1 || compLkRespLoc_firstReqAbt));
  assign _zz_8 = ({63'd0,1'b1} <<< compLkRespLoc_rCurTxnId);
  assign io_lkRespLoc_ready = (compLkRespLoc_stateReg == compLkRespLoc_enumDef_WAIT_RESP);
  assign io_axi_ar_payload_addr = {36'd0, _zz_io_axi_ar_payload_addr};
  assign io_axi_ar_payload_id = compLkRespLoc_rLkResp_payload_txnId;
  assign io_axi_ar_payload_len = (_zz_io_axi_ar_payload_len - 8'h01);
  assign io_axi_ar_payload_size = 3'b110;
  assign io_axi_ar_payload_burst = 2'b01;
  assign io_axi_ar_valid = (compLkRespLoc_stateReg == compLkRespLoc_enumDef_LOCAL_RD_REQ);
  assign compLkRespRmt_wantExit = 1'b0;
  always @(*) begin
    compLkRespRmt_wantStart = 1'b0;
    case(compLkRespRmt_stateReg)
      compLkRespRmt_enumDef_WAIT_RESP : begin
      end
      compLkRespRmt_enumDef_RMT_RD_CONSUME : begin
      end
      default : begin
        compLkRespRmt_wantStart = 1'b1;
      end
    endcase
  end

  assign compLkRespRmt_wantKill = 1'b0;
  assign io_lkRespRmt_fire = (io_lkRespRmt_valid && io_lkRespRmt_ready);
  assign compLkRespRmt_txnOffs = ({6'd0,io_lkRespRmt_payload_txnId} <<< 6);
  assign io_lkRespRmt_fire_1 = (io_lkRespRmt_valid && io_lkRespRmt_ready);
  assign compLkRespRmt_getAllRlse = ((_zz_compLkRespRmt_getAllRlse == _zz_compLkRespRmt_getAllRlse_1) && (_zz_compLkRespRmt_getAllRlse_2 == _zz_compLkRespRmt_getAllRlse_3));
  assign compLkRespRmt_getAllLkResp = ((_zz_compLkRespRmt_getAllLkResp == _zz_compLkRespRmt_getAllLkResp_1) && (_zz_compLkRespRmt_getAllLkResp_2 == _zz_compLkRespRmt_getAllLkResp_3));
  assign _zz_cntRlseRespRmt_0 = _zz__zz_cntRlseRespRmt_0;
  assign _zz_9 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign _zz_cntLkHoldRmt_0 = _zz__zz_cntLkHoldRmt_0;
  assign _zz_10 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign _zz_cntLkWaitRmt_0 = _zz__zz_cntLkWaitRmt_0;
  assign _zz_11 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign compLkRespRmt_getAllRlseTimeOut = ((_zz_compLkRespRmt_getAllRlseTimeOut == _zz_compLkRespRmt_getAllRlseTimeOut_1) && (_zz_cntRlseRespRmt_0 == _zz_compLkRespRmt_getAllRlseTimeOut_4));
  assign when_TxnManCS_l261 = _zz_when_TxnManCS_l261;
  assign io_lkReqLoc_fire_1 = (io_lkReqLoc_valid && io_lkReqLoc_ready);
  assign io_lkReqRmt_fire_1 = (io_lkReqRmt_valid && io_lkReqRmt_ready);
  assign compLkRespRmt_firstReqAbt = ((when_TxnManCS_l261 && (! (io_lkReqLoc_fire_1 && (io_lkReqLoc_payload_txnId == compLkRespRmt_rCurTxnId)))) && (! (io_lkReqRmt_fire_1 && (io_lkReqRmt_payload_txnId == compLkRespRmt_rCurTxnId))));
  assign io_lkRespRmt_fire_2 = (io_lkRespRmt_valid && io_lkRespRmt_ready);
  assign when_TxnManCS_l259 = ((compLkRespRmt_rFire && ((compLkRespRmt_getAllRlse && compLkRespRmt_getAllLkResp) || (_zz_when_TxnManCS_l259 && compLkRespRmt_getAllRlseTimeOut))) && (_zz_when_TxnManCS_l259_1 || compLkRespRmt_firstReqAbt));
  assign _zz_12 = ({63'd0,1'b1} <<< compLkRespRmt_rCurTxnId);
  assign io_lkRespRmt_ready = (compLkRespRmt_stateReg == compLkRespRmt_enumDef_WAIT_RESP);
  assign io_rdRmt_ready = (compLkRespRmt_stateReg == compLkRespRmt_enumDef_RMT_RD_CONSUME);
  assign io_axi_r_ready = 1'b1;
  assign io_axi_b_ready = 1'b1;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  assign _zz_13 = ({63'd0,1'b1} <<< compAxiResp_rAxiBId);
  assign _zz_cntCmtRespLoc_0 = (_zz__zz_cntCmtRespLoc_0 + 6'h01);
  assign compTxnCmtLoc_wantExit = 1'b0;
  always @(*) begin
    compTxnCmtLoc_wantStart = 1'b0;
    case(compTxnCmtLoc_stateReg)
      compTxnCmtLoc_enumDef_CS_TXN : begin
      end
      compTxnCmtLoc_enumDef_LOCAL_AW : begin
      end
      compTxnCmtLoc_enumDef_LOCAL_W : begin
      end
      default : begin
        compTxnCmtLoc_wantStart = 1'b1;
      end
    endcase
  end

  assign compTxnCmtLoc_wantKill = 1'b0;
  assign compTxnCmtLoc_txnOffs = ({6'd0,compTxnCmtLoc_curTxnId} <<< 6);
  assign _zz_cntCmtReqLoc_0 = _zz__zz_cntCmtReqLoc_0;
  assign _zz_14 = ({63'd0,1'b1} <<< compTxnCmtLoc_curTxnId);
  assign _zz_compTxnCmtLoc_cmtTxn_nId = (compTxnCmtLoc_txnOffs + _zz__zz_compTxnCmtLoc_cmtTxn_nId);
  assign _zz_compTxnCmtLoc_cmtTxn_nId_1 = _zz_txnWrMemLoc_port0;
  assign compTxnCmtLoc_cmtTxn_nId = _zz_compTxnCmtLoc_cmtTxn_nId_1[0 : 0];
  assign compTxnCmtLoc_cmtTxn_tId = _zz_compTxnCmtLoc_cmtTxn_nId_1[22 : 1];
  assign compTxnCmtLoc_cmtTxn_tabId = _zz_compTxnCmtLoc_cmtTxn_nId_1[25 : 23];
  assign _zz_compTxnCmtLoc_cmtTxn_lkType = _zz_compTxnCmtLoc_cmtTxn_nId_1[27 : 26];
  assign compTxnCmtLoc_cmtTxn_lkType = _zz_compTxnCmtLoc_cmtTxn_lkType;
  assign compTxnCmtLoc_cmtTxn_wLen = _zz_compTxnCmtLoc_cmtTxn_nId_1[30 : 28];
  assign compTxnCmtLoc_getAllLkResp = ((_zz_compTxnCmtLoc_getAllLkResp == _zz_compTxnCmtLoc_getAllLkResp_1) && (_zz_compTxnCmtLoc_getAllLkResp_2 == _zz_compTxnCmtLoc_getAllLkResp_3));
  assign io_axi_aw_payload_addr = {36'd0, _zz_io_axi_aw_payload_addr};
  assign io_axi_aw_payload_id = compTxnCmtLoc_curTxnId;
  assign io_axi_aw_payload_len = (_zz_io_axi_aw_payload_len - 8'h01);
  assign io_axi_aw_payload_size = 3'b110;
  assign io_axi_aw_payload_burst = 2'b01;
  assign io_axi_aw_valid = (compTxnCmtLoc_stateReg == compTxnCmtLoc_enumDef_LOCAL_AW);
  assign io_axi_w_payload_data = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
  assign io_axi_w_payload_last = (compTxnCmtLoc_nBeat == _zz_io_axi_w_payload_last);
  assign io_axi_w_valid = (compTxnCmtLoc_stateReg == compTxnCmtLoc_enumDef_LOCAL_W);
  assign compLkRlseLoc_wantExit = 1'b0;
  always @(*) begin
    compLkRlseLoc_wantStart = 1'b0;
    case(compLkRlseLoc_stateReg)
      compLkRlseLoc_enumDef_CS_TXN : begin
      end
      compLkRlseLoc_enumDef_LK_RLSE : begin
      end
      default : begin
        compLkRlseLoc_wantStart = 1'b1;
      end
    endcase
  end

  assign compLkRlseLoc_wantKill = 1'b0;
  assign compLkRlseLoc_txnOffs = ({6'd0,compLkRlseLoc_curTxnId} <<< 6);
  assign _zz_cntRlseReqLoc_0 = _zz__zz_cntRlseReqLoc_0;
  assign _zz_15 = ({63'd0,1'b1} <<< compLkRlseLoc_curTxnId);
  assign _zz_compLkRlseLoc_lkItem_nId = (compLkRlseLoc_txnOffs + _zz__zz_compLkRlseLoc_lkItem_nId);
  assign _zz_compLkRlseLoc_lkItem_nId_1 = _zz_lkMemLoc_port0;
  assign compLkRlseLoc_lkItem_nId = _zz_compLkRlseLoc_lkItem_nId_1[0 : 0];
  assign compLkRlseLoc_lkItem_tId = _zz_compLkRlseLoc_lkItem_nId_1[22 : 1];
  assign compLkRlseLoc_lkItem_tabId = _zz_compLkRlseLoc_lkItem_nId_1[25 : 23];
  assign compLkRlseLoc_lkItem_snId = _zz_compLkRlseLoc_lkItem_nId_1[26 : 26];
  assign compLkRlseLoc_lkItem_txnId = _zz_compLkRlseLoc_lkItem_nId_1[32 : 27];
  assign _zz_compLkRlseLoc_lkItem_lkType = _zz_compLkRlseLoc_lkItem_nId_1[34 : 33];
  assign compLkRlseLoc_lkItem_lkType = _zz_compLkRlseLoc_lkItem_lkType;
  assign compLkRlseLoc_lkItem_lkRelease = _zz_compLkRlseLoc_lkItem_nId_1[35];
  assign compLkRlseLoc_lkItem_txnAbt = _zz_compLkRlseLoc_lkItem_nId_1[36];
  assign compLkRlseLoc_lkItem_lkIdx = _zz_compLkRlseLoc_lkItem_nId_1[42 : 37];
  assign compLkRlseLoc_lkItem_wLen = _zz_compLkRlseLoc_lkItem_nId_1[45 : 43];
  assign _zz_compLkRlseLoc_lkItem_respType = _zz_compLkRlseLoc_lkItem_nId_1[47 : 46];
  assign compLkRlseLoc_lkItem_respType = _zz_compLkRlseLoc_lkItem_respType;
  assign compLkRlseLoc_lkItem_lkWaited = _zz_compLkRlseLoc_lkItem_nId_1[48];
  assign compLkRlseLoc_getAllLkResp = ((_zz_compLkRlseLoc_getAllLkResp == _zz_compLkRlseLoc_getAllLkResp_1) && (_zz_compLkRlseLoc_getAllLkResp_2 == _zz_compLkRlseLoc_getAllLkResp_3));
  assign _zz_lkReqRlseLoc_payload_txnAbt = _zz__zz_lkReqRlseLoc_payload_txnAbt;
  assign _zz_lkReqRlseLoc_payload_txnTimeOut = _zz__zz_lkReqRlseLoc_payload_txnTimeOut;
  assign _zz_lkReqRlseLoc_payload_lkType = compLkRlseLoc_lkItem_lkType;
  always @(*) begin
    _zz_lkReqRlseLoc_payload_lkRelease = compLkRlseLoc_lkItem_lkRelease;
    _zz_lkReqRlseLoc_payload_lkRelease = 1'b1;
  end

  always @(*) begin
    _zz_lkReqRlseLoc_payload_txnAbt_1 = compLkRlseLoc_lkItem_txnAbt;
    _zz_lkReqRlseLoc_payload_txnAbt_1 = _zz_lkReqRlseLoc_payload_txnAbt;
  end

  always @(*) begin
    _zz_lkReqRlseLoc_payload_lkIdx = compLkRlseLoc_lkItem_lkIdx;
    _zz_lkReqRlseLoc_payload_lkIdx = compLkRlseLoc_lkItem_lkIdx;
  end

  assign _zz_lkReqRlseLoc_payload_txnTimeOut_1 = _zz_lkReqRlseLoc_payload_txnTimeOut;
  assign lkReqRlseLoc_payload_nId = compLkRlseLoc_lkItem_nId;
  assign lkReqRlseLoc_payload_tId = compLkRlseLoc_lkItem_tId;
  assign lkReqRlseLoc_payload_tabId = compLkRlseLoc_lkItem_tabId;
  assign lkReqRlseLoc_payload_snId = compLkRlseLoc_lkItem_snId;
  assign lkReqRlseLoc_payload_txnId = compLkRlseLoc_lkItem_txnId;
  assign lkReqRlseLoc_payload_lkType = _zz_lkReqRlseLoc_payload_lkType;
  assign lkReqRlseLoc_payload_lkRelease = _zz_lkReqRlseLoc_payload_lkRelease;
  assign lkReqRlseLoc_payload_txnTimeOut = _zz_lkReqRlseLoc_payload_txnTimeOut_1;
  assign lkReqRlseLoc_payload_txnAbt = _zz_lkReqRlseLoc_payload_txnAbt_1;
  assign lkReqRlseLoc_payload_lkIdx = _zz_lkReqRlseLoc_payload_lkIdx;
  assign lkReqRlseLoc_payload_wLen = compLkRlseLoc_lkItem_wLen;
  assign compLkRlseRmt_wantExit = 1'b0;
  always @(*) begin
    compLkRlseRmt_wantStart = 1'b0;
    case(compLkRlseRmt_stateReg)
      compLkRlseRmt_enumDef_CS_TXN : begin
      end
      compLkRlseRmt_enumDef_RMT_LK_RLSE : begin
      end
      compLkRlseRmt_enumDef_RMT_WR : begin
      end
      default : begin
        compLkRlseRmt_wantStart = 1'b1;
      end
    endcase
  end

  assign compLkRlseRmt_wantKill = 1'b0;
  assign compLkRlseRmt_txnOffs = ({6'd0,compLkRlseRmt_curTxnId} <<< 6);
  assign _zz_cntRlseReqRmt_0 = _zz__zz_cntRlseReqRmt_0;
  assign _zz_16 = ({63'd0,1'b1} <<< compLkRlseRmt_curTxnId);
  assign _zz_17 = _zz_16[0];
  assign _zz_18 = _zz_16[1];
  assign _zz_19 = _zz_16[2];
  assign _zz_20 = _zz_16[3];
  assign _zz_21 = _zz_16[4];
  assign _zz_22 = _zz_16[5];
  assign _zz_23 = _zz_16[6];
  assign _zz_24 = _zz_16[7];
  assign _zz_25 = _zz_16[8];
  assign _zz_26 = _zz_16[9];
  assign _zz_27 = _zz_16[10];
  assign _zz_28 = _zz_16[11];
  assign _zz_29 = _zz_16[12];
  assign _zz_30 = _zz_16[13];
  assign _zz_31 = _zz_16[14];
  assign _zz_32 = _zz_16[15];
  assign _zz_33 = _zz_16[16];
  assign _zz_34 = _zz_16[17];
  assign _zz_35 = _zz_16[18];
  assign _zz_36 = _zz_16[19];
  assign _zz_37 = _zz_16[20];
  assign _zz_38 = _zz_16[21];
  assign _zz_39 = _zz_16[22];
  assign _zz_40 = _zz_16[23];
  assign _zz_41 = _zz_16[24];
  assign _zz_42 = _zz_16[25];
  assign _zz_43 = _zz_16[26];
  assign _zz_44 = _zz_16[27];
  assign _zz_45 = _zz_16[28];
  assign _zz_46 = _zz_16[29];
  assign _zz_47 = _zz_16[30];
  assign _zz_48 = _zz_16[31];
  assign _zz_49 = _zz_16[32];
  assign _zz_50 = _zz_16[33];
  assign _zz_51 = _zz_16[34];
  assign _zz_52 = _zz_16[35];
  assign _zz_53 = _zz_16[36];
  assign _zz_54 = _zz_16[37];
  assign _zz_55 = _zz_16[38];
  assign _zz_56 = _zz_16[39];
  assign _zz_57 = _zz_16[40];
  assign _zz_58 = _zz_16[41];
  assign _zz_59 = _zz_16[42];
  assign _zz_60 = _zz_16[43];
  assign _zz_61 = _zz_16[44];
  assign _zz_62 = _zz_16[45];
  assign _zz_63 = _zz_16[46];
  assign _zz_64 = _zz_16[47];
  assign _zz_65 = _zz_16[48];
  assign _zz_66 = _zz_16[49];
  assign _zz_67 = _zz_16[50];
  assign _zz_68 = _zz_16[51];
  assign _zz_69 = _zz_16[52];
  assign _zz_70 = _zz_16[53];
  assign _zz_71 = _zz_16[54];
  assign _zz_72 = _zz_16[55];
  assign _zz_73 = _zz_16[56];
  assign _zz_74 = _zz_16[57];
  assign _zz_75 = _zz_16[58];
  assign _zz_76 = _zz_16[59];
  assign _zz_77 = _zz_16[60];
  assign _zz_78 = _zz_16[61];
  assign _zz_79 = _zz_16[62];
  assign _zz_80 = _zz_16[63];
  assign _zz_compLkRlseRmt_lkItem_nId = (compLkRlseRmt_txnOffs + _zz__zz_compLkRlseRmt_lkItem_nId);
  assign _zz_compLkRlseRmt_lkItem_nId_1 = _zz_lkMemRmt_port0;
  assign compLkRlseRmt_lkItem_nId = _zz_compLkRlseRmt_lkItem_nId_1[0 : 0];
  assign compLkRlseRmt_lkItem_tId = _zz_compLkRlseRmt_lkItem_nId_1[22 : 1];
  assign compLkRlseRmt_lkItem_tabId = _zz_compLkRlseRmt_lkItem_nId_1[25 : 23];
  assign compLkRlseRmt_lkItem_snId = _zz_compLkRlseRmt_lkItem_nId_1[26 : 26];
  assign compLkRlseRmt_lkItem_txnId = _zz_compLkRlseRmt_lkItem_nId_1[32 : 27];
  assign _zz_compLkRlseRmt_lkItem_lkType = _zz_compLkRlseRmt_lkItem_nId_1[34 : 33];
  assign compLkRlseRmt_lkItem_lkType = _zz_compLkRlseRmt_lkItem_lkType;
  assign compLkRlseRmt_lkItem_lkRelease = _zz_compLkRlseRmt_lkItem_nId_1[35];
  assign compLkRlseRmt_lkItem_txnAbt = _zz_compLkRlseRmt_lkItem_nId_1[36];
  assign compLkRlseRmt_lkItem_lkIdx = _zz_compLkRlseRmt_lkItem_nId_1[42 : 37];
  assign compLkRlseRmt_lkItem_wLen = _zz_compLkRlseRmt_lkItem_nId_1[45 : 43];
  assign _zz_compLkRlseRmt_lkItem_respType = _zz_compLkRlseRmt_lkItem_nId_1[47 : 46];
  assign compLkRlseRmt_lkItem_respType = _zz_compLkRlseRmt_lkItem_respType;
  assign compLkRlseRmt_lkItem_lkWaited = _zz_compLkRlseRmt_lkItem_nId_1[48];
  assign compLkRlseRmt_getAllLkResp = ((_zz_compLkRlseRmt_getAllLkResp == _zz_compLkRlseRmt_getAllLkResp_1) && (_zz_compLkRlseRmt_getAllLkResp_2 == _zz_compLkRlseRmt_getAllLkResp_3));
  assign _zz_lkReqRlseRmt_payload_txnAbt = _zz__zz_lkReqRlseRmt_payload_txnAbt;
  assign _zz_lkReqRlseRmt_payload_txnTimeOut = _zz__zz_lkReqRlseRmt_payload_txnTimeOut;
  assign _zz_lkReqRlseRmt_payload_lkType = compLkRlseRmt_lkItem_lkType;
  always @(*) begin
    _zz_lkReqRlseRmt_payload_lkRelease = compLkRlseRmt_lkItem_lkRelease;
    _zz_lkReqRlseRmt_payload_lkRelease = 1'b1;
  end

  always @(*) begin
    _zz_lkReqRlseRmt_payload_txnAbt_1 = compLkRlseRmt_lkItem_txnAbt;
    _zz_lkReqRlseRmt_payload_txnAbt_1 = _zz_lkReqRlseRmt_payload_txnAbt;
  end

  always @(*) begin
    _zz_lkReqRlseRmt_payload_lkIdx = compLkRlseRmt_lkItem_lkIdx;
    _zz_lkReqRlseRmt_payload_lkIdx = compLkRlseRmt_lkItem_lkIdx;
  end

  assign _zz_lkReqRlseRmt_payload_txnTimeOut_1 = _zz_lkReqRlseRmt_payload_txnTimeOut;
  assign lkReqRlseRmt_payload_nId = compLkRlseRmt_lkItem_nId;
  assign lkReqRlseRmt_payload_tId = compLkRlseRmt_lkItem_tId;
  assign lkReqRlseRmt_payload_tabId = compLkRlseRmt_lkItem_tabId;
  assign lkReqRlseRmt_payload_snId = compLkRlseRmt_lkItem_snId;
  assign lkReqRlseRmt_payload_txnId = compLkRlseRmt_lkItem_txnId;
  assign lkReqRlseRmt_payload_lkType = _zz_lkReqRlseRmt_payload_lkType;
  assign lkReqRlseRmt_payload_lkRelease = _zz_lkReqRlseRmt_payload_lkRelease;
  assign lkReqRlseRmt_payload_txnTimeOut = _zz_lkReqRlseRmt_payload_txnTimeOut_1;
  assign lkReqRlseRmt_payload_txnAbt = _zz_lkReqRlseRmt_payload_txnAbt_1;
  assign lkReqRlseRmt_payload_lkIdx = _zz_lkReqRlseRmt_payload_lkIdx;
  assign lkReqRlseRmt_payload_wLen = compLkRlseRmt_lkItem_wLen;
  assign io_wrRmt_valid = (compLkRlseRmt_stateReg == compLkRlseRmt_enumDef_RMT_WR);
  assign io_wrRmt_payload = 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
  assign compTimeOut_wantExit = 1'b0;
  always @(*) begin
    compTimeOut_wantStart = 1'b0;
    case(compTimeOut_stateReg)
      compTimeOut_enumDef_IDLE : begin
      end
      compTimeOut_enumDef_COUNT : begin
      end
      default : begin
        compTimeOut_wantStart = 1'b1;
      end
    endcase
  end

  assign compTimeOut_wantKill = 1'b0;
  assign compLoadTxn_wantExit = 1'b0;
  always @(*) begin
    compLoadTxn_wantStart = 1'b0;
    case(compLoadTxn_stateReg)
      compLoadTxn_enumDef_IDLE : begin
      end
      compLoadTxn_enumDef_CS_TXN : begin
      end
      compLoadTxn_enumDef_RD_CMDAXI : begin
      end
      compLoadTxn_enumDef_LD_TXN : begin
      end
      default : begin
        compLoadTxn_wantStart = 1'b1;
      end
    endcase
  end

  assign compLoadTxn_wantKill = 1'b0;
  assign compLoadTxn_txnOffs = ({6'd0,compLoadTxn_curTxnId} <<< 6);
  assign io_cmdAxi_ar_payload_addr = {23'd0, _zz_io_cmdAxi_ar_payload_addr};
  assign io_cmdAxi_ar_payload_id = 6'h0;
  assign io_cmdAxi_ar_payload_len = {4'd0, _zz_io_cmdAxi_ar_payload_len};
  assign io_cmdAxi_ar_payload_size = 3'b110;
  assign io_cmdAxi_ar_payload_burst = 2'b01;
  assign io_cmdAxi_r_fire = (io_cmdAxi_r_valid && io_cmdAxi_r_ready);
  assign io_cmdAxi_r_fire_1 = (io_cmdAxi_r_valid && io_cmdAxi_r_ready);
  assign compLoadTxn_cmdAxiDataSlice_0 = compLoadTxn_rCmdAxiData[63 : 0];
  assign compLoadTxn_cmdAxiDataSlice_1 = compLoadTxn_rCmdAxiData[127 : 64];
  assign compLoadTxn_cmdAxiDataSlice_2 = compLoadTxn_rCmdAxiData[191 : 128];
  assign compLoadTxn_cmdAxiDataSlice_3 = compLoadTxn_rCmdAxiData[255 : 192];
  assign compLoadTxn_cmdAxiDataSlice_4 = compLoadTxn_rCmdAxiData[319 : 256];
  assign compLoadTxn_cmdAxiDataSlice_5 = compLoadTxn_rCmdAxiData[383 : 320];
  assign compLoadTxn_cmdAxiDataSlice_6 = compLoadTxn_rCmdAxiData[447 : 384];
  assign compLoadTxn_cmdAxiDataSlice_7 = compLoadTxn_rCmdAxiData[511 : 448];
  always @(*) begin
    compLoadTxn_cntTxnWordInLine_willIncrement = 1'b0;
    if(compLoadTxn_rTxnMemLd) begin
      compLoadTxn_cntTxnWordInLine_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    compLoadTxn_cntTxnWordInLine_willClear = 1'b0;
    case(compLoadTxn_stateReg)
      compLoadTxn_enumDef_IDLE : begin
      end
      compLoadTxn_enumDef_CS_TXN : begin
      end
      compLoadTxn_enumDef_RD_CMDAXI : begin
        if(io_cmdAxi_ar_fire) begin
          compLoadTxn_cntTxnWordInLine_willClear = 1'b1;
        end
      end
      compLoadTxn_enumDef_LD_TXN : begin
      end
      default : begin
      end
    endcase
  end

  assign compLoadTxn_cntTxnWordInLine_willOverflowIfInc = (compLoadTxn_cntTxnWordInLine_value == 3'b111);
  assign compLoadTxn_cntTxnWordInLine_willOverflow = (compLoadTxn_cntTxnWordInLine_willOverflowIfInc && compLoadTxn_cntTxnWordInLine_willIncrement);
  always @(*) begin
    compLoadTxn_cntTxnWordInLine_valueNext = (compLoadTxn_cntTxnWordInLine_value + _zz_compLoadTxn_cntTxnWordInLine_valueNext);
    if(compLoadTxn_cntTxnWordInLine_willClear) begin
      compLoadTxn_cntTxnWordInLine_valueNext = 3'b000;
    end
  end

  always @(*) begin
    compLoadTxn_cntTxnWord_willIncrement = 1'b0;
    if(compLoadTxn_rTxnMemLd) begin
      compLoadTxn_cntTxnWord_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    compLoadTxn_cntTxnWord_willClear = 1'b0;
    case(compLoadTxn_stateReg)
      compLoadTxn_enumDef_IDLE : begin
      end
      compLoadTxn_enumDef_CS_TXN : begin
      end
      compLoadTxn_enumDef_RD_CMDAXI : begin
        if(io_cmdAxi_ar_fire) begin
          compLoadTxn_cntTxnWord_willClear = 1'b1;
        end
      end
      compLoadTxn_enumDef_LD_TXN : begin
      end
      default : begin
      end
    endcase
  end

  assign compLoadTxn_cntTxnWord_willOverflowIfInc = (compLoadTxn_cntTxnWord_value == 6'h3f);
  assign compLoadTxn_cntTxnWord_willOverflow = (compLoadTxn_cntTxnWord_willOverflowIfInc && compLoadTxn_cntTxnWord_willIncrement);
  always @(*) begin
    compLoadTxn_cntTxnWord_valueNext = (compLoadTxn_cntTxnWord_value + _zz_compLoadTxn_cntTxnWord_valueNext);
    if(compLoadTxn_cntTxnWord_willClear) begin
      compLoadTxn_cntTxnWord_valueNext = 6'h0;
    end
  end

  assign compLoadTxn_bitsBuff = _zz_compLoadTxn_bitsBuff;
  assign compLoadTxn_txnBuff = {{{{compLoadTxn_bitsBuff[0 : 0],compLoadTxn_bitsBuff[39 : 18]},compLoadTxn_bitsBuff[14 : 12]},compLoadTxn_bitsBuff[43 : 42]},compLoadTxn_bitsBuff[48 : 46]};
  assign io_cmdAxi_ar_valid = (compLoadTxn_stateReg == compLoadTxn_enumDef_RD_CMDAXI);
  assign io_cmdAxi_r_ready = ((((compLoadTxn_stateReg == compLoadTxn_enumDef_LD_TXN) && (compLoadTxn_cntTxnWordInLine_value == 3'b000)) && (! compLoadTxn_rCmdAxiFire)) ? 1'b1 : 1'b0);
  assign when_TxnManCS_l672 = ((((((((((((((_zz_when_TxnManCS_l672 && rRlseDone_52) && rRlseDone_53) && rRlseDone_54) && rRlseDone_55) && rRlseDone_56) && rRlseDone_57) && rRlseDone_58) && rRlseDone_59) && rRlseDone_60) && rRlseDone_61) && rRlseDone_62) && rRlseDone_63) && (io_cntTxnLd == io_txnNumTotal)) && (! io_done));
  assign clkCnt_wantExit = 1'b0;
  always @(*) begin
    clkCnt_wantStart = 1'b0;
    case(clkCnt_stateReg)
      clkCnt_enumDef_IDLE : begin
      end
      clkCnt_enumDef_CNT : begin
      end
      default : begin
        clkCnt_wantStart = 1'b1;
      end
    endcase
  end

  assign clkCnt_wantKill = 1'b0;
  always @(*) begin
    compLkReq_stateNext = compLkReq_stateReg;
    case(compLkReq_stateReg)
      compLkReq_enumDef_CS_TXN : begin
        if(compLkReq_txnMemRd_fire) begin
          compLkReq_stateNext = compLkReq_enumDef_RD_TXN;
        end
      end
      compLkReq_enumDef_RD_TXN : begin
        if(when_TxnManCS_l128) begin
          compLkReq_stateNext = compLkReq_enumDef_CS_TXN;
        end
      end
      default : begin
      end
    endcase
    if(compLkReq_wantStart) begin
      compLkReq_stateNext = compLkReq_enumDef_CS_TXN;
    end
    if(compLkReq_wantKill) begin
      compLkReq_stateNext = compLkReq_enumDef_BOOT;
    end
  end

  assign compLkReq_txnMemRd_fire = (compLkReq_txnMemRd_valid && compLkReq_txnMemRd_ready);
  assign _zz_compLkReq_txnMemRdCmd_payload = (_zz__zz_compLkReq_txnMemRdCmd_payload + 12'h001);
  assign _zz_82 = ({63'd0,1'b1} <<< compLkReq_curTxnId);
  assign _zz_cntLkReqLoc_0 = (_zz__zz_cntLkReqLoc_0 + 6'h01);
  assign _zz_83 = ({63'd0,1'b1} <<< compLkReq_curTxnId);
  assign _zz_cntLkReqRmt_0 = (_zz__zz_cntLkReqRmt_0 + 6'h01);
  assign when_TxnManCS_l106 = ((compLkReq_txnMemRd_payload_lkType == LkT_wr) || (compLkReq_txnMemRd_payload_lkType == LkT_raw));
  assign _zz_cntLkReqWrLoc_0 = _zz__zz_cntLkReqWrLoc_0;
  assign _zz_84 = ({63'd0,1'b1} <<< compLkReq_curTxnId);
  assign _zz_cntLkReqWrLoc_0_1 = (_zz_cntLkReqWrLoc_0 + 6'h01);
  assign _zz_cntLkReqWrRmt_0 = _zz__zz_cntLkReqWrRmt_0;
  assign _zz_85 = ({63'd0,1'b1} <<< compLkReq_curTxnId);
  assign _zz_cntLkReqWrRmt_0_1 = (_zz_cntLkReqWrRmt_0 + 6'h01);
  assign when_TxnManCS_l128 = ((compLkReq_lkReqFire && (compLkReq_reqIdx == _zz_when_TxnManCS_l128)) || _zz_when_TxnManCS_l128_1);
  assign _zz_86 = ({63'd0,1'b1} <<< compLkReq_curTxnId);
  always @(*) begin
    compLkRespLoc_stateNext = compLkRespLoc_stateReg;
    case(compLkRespLoc_stateReg)
      compLkRespLoc_enumDef_WAIT_RESP : begin
        if(io_lkRespLoc_fire_3) begin
          case(io_lkRespLoc_payload_respType)
            LockRespType_grant : begin
              case(io_lkRespLoc_payload_lkType)
                LkT_rd : begin
                  compLkRespLoc_stateNext = compLkRespLoc_enumDef_LOCAL_RD_REQ;
                end
                LkT_wr : begin
                end
                LkT_raw : begin
                  compLkRespLoc_stateNext = compLkRespLoc_enumDef_LOCAL_RD_REQ;
                end
                default : begin
                end
              endcase
            end
            LockRespType_waiting : begin
            end
            LockRespType_abort : begin
            end
            default : begin
            end
          endcase
        end
      end
      compLkRespLoc_enumDef_LOCAL_RD_REQ : begin
        if(io_axi_ar_fire) begin
          compLkRespLoc_stateNext = compLkRespLoc_enumDef_WAIT_RESP;
        end
      end
      default : begin
      end
    endcase
    if(compLkRespLoc_wantStart) begin
      compLkRespLoc_stateNext = compLkRespLoc_enumDef_WAIT_RESP;
    end
    if(compLkRespLoc_wantKill) begin
      compLkRespLoc_stateNext = compLkRespLoc_enumDef_BOOT;
    end
  end

  assign io_lkRespLoc_fire_3 = (io_lkRespLoc_valid && io_lkRespLoc_ready);
  assign _zz_cntLkRespLoc_0 = _zz__zz_cntLkRespLoc_0;
  assign _zz_87 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign _zz_88 = _zz_87[0];
  assign _zz_89 = _zz_87[1];
  assign _zz_90 = _zz_87[2];
  assign _zz_91 = _zz_87[3];
  assign _zz_92 = _zz_87[4];
  assign _zz_93 = _zz_87[5];
  assign _zz_94 = _zz_87[6];
  assign _zz_95 = _zz_87[7];
  assign _zz_96 = _zz_87[8];
  assign _zz_97 = _zz_87[9];
  assign _zz_98 = _zz_87[10];
  assign _zz_99 = _zz_87[11];
  assign _zz_100 = _zz_87[12];
  assign _zz_101 = _zz_87[13];
  assign _zz_102 = _zz_87[14];
  assign _zz_103 = _zz_87[15];
  assign _zz_104 = _zz_87[16];
  assign _zz_105 = _zz_87[17];
  assign _zz_106 = _zz_87[18];
  assign _zz_107 = _zz_87[19];
  assign _zz_108 = _zz_87[20];
  assign _zz_109 = _zz_87[21];
  assign _zz_110 = _zz_87[22];
  assign _zz_111 = _zz_87[23];
  assign _zz_112 = _zz_87[24];
  assign _zz_113 = _zz_87[25];
  assign _zz_114 = _zz_87[26];
  assign _zz_115 = _zz_87[27];
  assign _zz_116 = _zz_87[28];
  assign _zz_117 = _zz_87[29];
  assign _zz_118 = _zz_87[30];
  assign _zz_119 = _zz_87[31];
  assign _zz_120 = _zz_87[32];
  assign _zz_121 = _zz_87[33];
  assign _zz_122 = _zz_87[34];
  assign _zz_123 = _zz_87[35];
  assign _zz_124 = _zz_87[36];
  assign _zz_125 = _zz_87[37];
  assign _zz_126 = _zz_87[38];
  assign _zz_127 = _zz_87[39];
  assign _zz_128 = _zz_87[40];
  assign _zz_129 = _zz_87[41];
  assign _zz_130 = _zz_87[42];
  assign _zz_131 = _zz_87[43];
  assign _zz_132 = _zz_87[44];
  assign _zz_133 = _zz_87[45];
  assign _zz_134 = _zz_87[46];
  assign _zz_135 = _zz_87[47];
  assign _zz_136 = _zz_87[48];
  assign _zz_137 = _zz_87[49];
  assign _zz_138 = _zz_87[50];
  assign _zz_139 = _zz_87[51];
  assign _zz_140 = _zz_87[52];
  assign _zz_141 = _zz_87[53];
  assign _zz_142 = _zz_87[54];
  assign _zz_143 = _zz_87[55];
  assign _zz_144 = _zz_87[56];
  assign _zz_145 = _zz_87[57];
  assign _zz_146 = _zz_87[58];
  assign _zz_147 = _zz_87[59];
  assign _zz_148 = _zz_87[60];
  assign _zz_149 = _zz_87[61];
  assign _zz_150 = _zz_87[62];
  assign _zz_151 = _zz_87[63];
  assign _zz_cntLkRespLoc_0_1 = (_zz_cntLkRespLoc_0 + 6'h01);
  assign when_TxnManCS_l179 = (io_lkRespLoc_payload_lkType != LkT_insTab);
  assign _zz_cntLkHoldLoc_0_1 = (_zz_cntLkHoldLoc_0 + 6'h01);
  assign _zz_cntLkHoldWrLoc_0 = _zz__zz_cntLkHoldWrLoc_0;
  assign _zz_152 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign _zz_153 = _zz_152[0];
  assign _zz_154 = _zz_152[1];
  assign _zz_155 = _zz_152[2];
  assign _zz_156 = _zz_152[3];
  assign _zz_157 = _zz_152[4];
  assign _zz_158 = _zz_152[5];
  assign _zz_159 = _zz_152[6];
  assign _zz_160 = _zz_152[7];
  assign _zz_161 = _zz_152[8];
  assign _zz_162 = _zz_152[9];
  assign _zz_163 = _zz_152[10];
  assign _zz_164 = _zz_152[11];
  assign _zz_165 = _zz_152[12];
  assign _zz_166 = _zz_152[13];
  assign _zz_167 = _zz_152[14];
  assign _zz_168 = _zz_152[15];
  assign _zz_169 = _zz_152[16];
  assign _zz_170 = _zz_152[17];
  assign _zz_171 = _zz_152[18];
  assign _zz_172 = _zz_152[19];
  assign _zz_173 = _zz_152[20];
  assign _zz_174 = _zz_152[21];
  assign _zz_175 = _zz_152[22];
  assign _zz_176 = _zz_152[23];
  assign _zz_177 = _zz_152[24];
  assign _zz_178 = _zz_152[25];
  assign _zz_179 = _zz_152[26];
  assign _zz_180 = _zz_152[27];
  assign _zz_181 = _zz_152[28];
  assign _zz_182 = _zz_152[29];
  assign _zz_183 = _zz_152[30];
  assign _zz_184 = _zz_152[31];
  assign _zz_185 = _zz_152[32];
  assign _zz_186 = _zz_152[33];
  assign _zz_187 = _zz_152[34];
  assign _zz_188 = _zz_152[35];
  assign _zz_189 = _zz_152[36];
  assign _zz_190 = _zz_152[37];
  assign _zz_191 = _zz_152[38];
  assign _zz_192 = _zz_152[39];
  assign _zz_193 = _zz_152[40];
  assign _zz_194 = _zz_152[41];
  assign _zz_195 = _zz_152[42];
  assign _zz_196 = _zz_152[43];
  assign _zz_197 = _zz_152[44];
  assign _zz_198 = _zz_152[45];
  assign _zz_199 = _zz_152[46];
  assign _zz_200 = _zz_152[47];
  assign _zz_201 = _zz_152[48];
  assign _zz_202 = _zz_152[49];
  assign _zz_203 = _zz_152[50];
  assign _zz_204 = _zz_152[51];
  assign _zz_205 = _zz_152[52];
  assign _zz_206 = _zz_152[53];
  assign _zz_207 = _zz_152[54];
  assign _zz_208 = _zz_152[55];
  assign _zz_209 = _zz_152[56];
  assign _zz_210 = _zz_152[57];
  assign _zz_211 = _zz_152[58];
  assign _zz_212 = _zz_152[59];
  assign _zz_213 = _zz_152[60];
  assign _zz_214 = _zz_152[61];
  assign _zz_215 = _zz_152[62];
  assign _zz_216 = _zz_152[63];
  assign _zz_cntLkHoldWrLoc_0_1 = (_zz_cntLkHoldWrLoc_0 + 6'h01);
  assign _zz_cntLkHoldWrLoc_0_2 = (_zz_cntLkHoldWrLoc_0 + 6'h01);
  assign _zz_cntLkWaitLoc_0_1 = (_zz_cntLkWaitLoc_0 + 6'h01);
  assign _zz_217 = ({63'd0,1'b1} <<< io_lkRespLoc_payload_txnId);
  assign _zz_cntLkRespLoc_0_2 = (_zz_cntLkRespLoc_0 + 6'h01);
  assign _zz_cntRlseRespLoc_0_1 = (_zz_cntRlseRespLoc_0 + 6'h01);
  assign when_TxnManCS_l214 = (((io_lkRespLoc_payload_respType == LockRespType_grant) && (! io_lkRespLoc_payload_lkWaited)) || (io_lkRespLoc_payload_respType == LockRespType_waiting));
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  always @(*) begin
    compLkRespRmt_stateNext = compLkRespRmt_stateReg;
    case(compLkRespRmt_stateReg)
      compLkRespRmt_enumDef_WAIT_RESP : begin
        if(io_lkRespRmt_fire_3) begin
          case(io_lkRespRmt_payload_respType)
            LockRespType_grant : begin
              case(io_lkRespRmt_payload_lkType)
                LkT_rd : begin
                  compLkRespRmt_stateNext = compLkRespRmt_enumDef_RMT_RD_CONSUME;
                end
                LkT_wr : begin
                end
                LkT_raw : begin
                  compLkRespRmt_stateNext = compLkRespRmt_enumDef_RMT_RD_CONSUME;
                end
                default : begin
                end
              endcase
            end
            LockRespType_waiting : begin
            end
            LockRespType_abort : begin
            end
            default : begin
            end
          endcase
        end
      end
      compLkRespRmt_enumDef_RMT_RD_CONSUME : begin
        if(io_rdRmt_fire) begin
          if(when_TxnManCS_l315) begin
            compLkRespRmt_stateNext = compLkRespRmt_enumDef_WAIT_RESP;
          end
        end
      end
      default : begin
      end
    endcase
    if(compLkRespRmt_wantStart) begin
      compLkRespRmt_stateNext = compLkRespRmt_enumDef_WAIT_RESP;
    end
    if(compLkRespRmt_wantKill) begin
      compLkRespRmt_stateNext = compLkRespRmt_enumDef_BOOT;
    end
  end

  assign io_lkRespRmt_fire_3 = (io_lkRespRmt_valid && io_lkRespRmt_ready);
  assign _zz_cntLkRespRmt_0 = _zz__zz_cntLkRespRmt_0;
  assign _zz_218 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign _zz_219 = _zz_218[0];
  assign _zz_220 = _zz_218[1];
  assign _zz_221 = _zz_218[2];
  assign _zz_222 = _zz_218[3];
  assign _zz_223 = _zz_218[4];
  assign _zz_224 = _zz_218[5];
  assign _zz_225 = _zz_218[6];
  assign _zz_226 = _zz_218[7];
  assign _zz_227 = _zz_218[8];
  assign _zz_228 = _zz_218[9];
  assign _zz_229 = _zz_218[10];
  assign _zz_230 = _zz_218[11];
  assign _zz_231 = _zz_218[12];
  assign _zz_232 = _zz_218[13];
  assign _zz_233 = _zz_218[14];
  assign _zz_234 = _zz_218[15];
  assign _zz_235 = _zz_218[16];
  assign _zz_236 = _zz_218[17];
  assign _zz_237 = _zz_218[18];
  assign _zz_238 = _zz_218[19];
  assign _zz_239 = _zz_218[20];
  assign _zz_240 = _zz_218[21];
  assign _zz_241 = _zz_218[22];
  assign _zz_242 = _zz_218[23];
  assign _zz_243 = _zz_218[24];
  assign _zz_244 = _zz_218[25];
  assign _zz_245 = _zz_218[26];
  assign _zz_246 = _zz_218[27];
  assign _zz_247 = _zz_218[28];
  assign _zz_248 = _zz_218[29];
  assign _zz_249 = _zz_218[30];
  assign _zz_250 = _zz_218[31];
  assign _zz_251 = _zz_218[32];
  assign _zz_252 = _zz_218[33];
  assign _zz_253 = _zz_218[34];
  assign _zz_254 = _zz_218[35];
  assign _zz_255 = _zz_218[36];
  assign _zz_256 = _zz_218[37];
  assign _zz_257 = _zz_218[38];
  assign _zz_258 = _zz_218[39];
  assign _zz_259 = _zz_218[40];
  assign _zz_260 = _zz_218[41];
  assign _zz_261 = _zz_218[42];
  assign _zz_262 = _zz_218[43];
  assign _zz_263 = _zz_218[44];
  assign _zz_264 = _zz_218[45];
  assign _zz_265 = _zz_218[46];
  assign _zz_266 = _zz_218[47];
  assign _zz_267 = _zz_218[48];
  assign _zz_268 = _zz_218[49];
  assign _zz_269 = _zz_218[50];
  assign _zz_270 = _zz_218[51];
  assign _zz_271 = _zz_218[52];
  assign _zz_272 = _zz_218[53];
  assign _zz_273 = _zz_218[54];
  assign _zz_274 = _zz_218[55];
  assign _zz_275 = _zz_218[56];
  assign _zz_276 = _zz_218[57];
  assign _zz_277 = _zz_218[58];
  assign _zz_278 = _zz_218[59];
  assign _zz_279 = _zz_218[60];
  assign _zz_280 = _zz_218[61];
  assign _zz_281 = _zz_218[62];
  assign _zz_282 = _zz_218[63];
  assign _zz_cntLkRespRmt_0_1 = (_zz_cntLkRespRmt_0 + 6'h01);
  assign when_TxnManCS_l272 = (io_lkRespRmt_payload_lkType != LkT_insTab);
  assign _zz_cntLkHoldRmt_0_1 = (_zz_cntLkHoldRmt_0 + 6'h01);
  assign _zz_cntLkHoldWrRmt_0 = _zz__zz_cntLkHoldWrRmt_0;
  assign _zz_283 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign _zz_284 = _zz_283[0];
  assign _zz_285 = _zz_283[1];
  assign _zz_286 = _zz_283[2];
  assign _zz_287 = _zz_283[3];
  assign _zz_288 = _zz_283[4];
  assign _zz_289 = _zz_283[5];
  assign _zz_290 = _zz_283[6];
  assign _zz_291 = _zz_283[7];
  assign _zz_292 = _zz_283[8];
  assign _zz_293 = _zz_283[9];
  assign _zz_294 = _zz_283[10];
  assign _zz_295 = _zz_283[11];
  assign _zz_296 = _zz_283[12];
  assign _zz_297 = _zz_283[13];
  assign _zz_298 = _zz_283[14];
  assign _zz_299 = _zz_283[15];
  assign _zz_300 = _zz_283[16];
  assign _zz_301 = _zz_283[17];
  assign _zz_302 = _zz_283[18];
  assign _zz_303 = _zz_283[19];
  assign _zz_304 = _zz_283[20];
  assign _zz_305 = _zz_283[21];
  assign _zz_306 = _zz_283[22];
  assign _zz_307 = _zz_283[23];
  assign _zz_308 = _zz_283[24];
  assign _zz_309 = _zz_283[25];
  assign _zz_310 = _zz_283[26];
  assign _zz_311 = _zz_283[27];
  assign _zz_312 = _zz_283[28];
  assign _zz_313 = _zz_283[29];
  assign _zz_314 = _zz_283[30];
  assign _zz_315 = _zz_283[31];
  assign _zz_316 = _zz_283[32];
  assign _zz_317 = _zz_283[33];
  assign _zz_318 = _zz_283[34];
  assign _zz_319 = _zz_283[35];
  assign _zz_320 = _zz_283[36];
  assign _zz_321 = _zz_283[37];
  assign _zz_322 = _zz_283[38];
  assign _zz_323 = _zz_283[39];
  assign _zz_324 = _zz_283[40];
  assign _zz_325 = _zz_283[41];
  assign _zz_326 = _zz_283[42];
  assign _zz_327 = _zz_283[43];
  assign _zz_328 = _zz_283[44];
  assign _zz_329 = _zz_283[45];
  assign _zz_330 = _zz_283[46];
  assign _zz_331 = _zz_283[47];
  assign _zz_332 = _zz_283[48];
  assign _zz_333 = _zz_283[49];
  assign _zz_334 = _zz_283[50];
  assign _zz_335 = _zz_283[51];
  assign _zz_336 = _zz_283[52];
  assign _zz_337 = _zz_283[53];
  assign _zz_338 = _zz_283[54];
  assign _zz_339 = _zz_283[55];
  assign _zz_340 = _zz_283[56];
  assign _zz_341 = _zz_283[57];
  assign _zz_342 = _zz_283[58];
  assign _zz_343 = _zz_283[59];
  assign _zz_344 = _zz_283[60];
  assign _zz_345 = _zz_283[61];
  assign _zz_346 = _zz_283[62];
  assign _zz_347 = _zz_283[63];
  assign _zz_cntLkHoldWrRmt_0_1 = (_zz_cntLkHoldWrRmt_0 + 6'h01);
  assign _zz_cntLkHoldWrRmt_0_2 = (_zz_cntLkHoldWrRmt_0 + 6'h01);
  assign _zz_cntLkWaitRmt_0_1 = (_zz_cntLkWaitRmt_0 + 6'h01);
  assign _zz_348 = ({63'd0,1'b1} <<< io_lkRespRmt_payload_txnId);
  assign _zz_cntLkRespRmt_0_2 = (_zz_cntLkRespRmt_0 + 6'h01);
  assign _zz_cntRlseRespRmt_0_1 = (_zz_cntRlseRespRmt_0 + 6'h01);
  assign when_TxnManCS_l303 = (((io_lkRespRmt_payload_respType == LockRespType_grant) && (! io_lkRespRmt_payload_lkWaited)) || (io_lkRespRmt_payload_respType == LockRespType_waiting));
  assign io_rdRmt_fire = (io_rdRmt_valid && io_rdRmt_ready);
  assign when_TxnManCS_l315 = (compLkRespRmt_nBeat == _zz_when_TxnManCS_l315);
  always @(*) begin
    compTxnCmtLoc_stateNext = compTxnCmtLoc_stateReg;
    case(compTxnCmtLoc_stateReg)
      compTxnCmtLoc_enumDef_CS_TXN : begin
        if(when_TxnManCS_l369) begin
          compTxnCmtLoc_stateNext = compTxnCmtLoc_enumDef_LOCAL_AW;
        end
      end
      compTxnCmtLoc_enumDef_LOCAL_AW : begin
        if(io_axi_aw_fire) begin
          compTxnCmtLoc_stateNext = compTxnCmtLoc_enumDef_LOCAL_W;
        end
      end
      compTxnCmtLoc_enumDef_LOCAL_W : begin
        if(io_axi_w_fire) begin
          if(io_axi_w_payload_last) begin
            compTxnCmtLoc_stateNext = compTxnCmtLoc_enumDef_CS_TXN;
          end
        end
      end
      default : begin
      end
    endcase
    if(compTxnCmtLoc_wantStart) begin
      compTxnCmtLoc_stateNext = compTxnCmtLoc_enumDef_CS_TXN;
    end
    if(compTxnCmtLoc_wantKill) begin
      compTxnCmtLoc_stateNext = compTxnCmtLoc_enumDef_BOOT;
    end
  end

  assign when_TxnManCS_l369 = (((compTxnCmtLoc_getAllLkResp && _zz_when_TxnManCS_l369) && (! _zz_when_TxnManCS_l369_1)) && (_zz_cntCmtReqLoc_0 < _zz_when_TxnManCS_l369_2));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign _zz_cntCmtReqLoc_0_1 = (_zz_cntCmtReqLoc_0 + 6'h01);
  always @(*) begin
    compLkRlseLoc_stateNext = compLkRlseLoc_stateReg;
    case(compLkRlseLoc_stateReg)
      compLkRlseLoc_enumDef_CS_TXN : begin
        if(when_TxnManCS_l440) begin
          compLkRlseLoc_stateNext = compLkRlseLoc_enumDef_LK_RLSE;
        end
      end
      compLkRlseLoc_enumDef_LK_RLSE : begin
        if(lkReqRlseLoc_fire) begin
          compLkRlseLoc_stateNext = compLkRlseLoc_enumDef_CS_TXN;
        end
      end
      default : begin
      end
    endcase
    if(compLkRlseLoc_wantStart) begin
      compLkRlseLoc_stateNext = compLkRlseLoc_enumDef_CS_TXN;
    end
    if(compLkRlseLoc_wantKill) begin
      compLkRlseLoc_stateNext = compLkRlseLoc_enumDef_BOOT;
    end
  end

  assign _zz_cntRlseReqWrLoc_0 = _zz__zz_cntRlseReqWrLoc_0;
  assign _zz_349 = ({63'd0,1'b1} <<< compLkRlseLoc_curTxnId);
  assign _zz_when_TxnManCS_l440 = _zz__zz_when_TxnManCS_l440;
  assign when_TxnManCS_l440 = ((((compLkRlseLoc_getAllLkResp && (_zz_lkReqRlseLoc_payload_txnAbt || _zz_when_TxnManCS_l440_1)) && ((_zz_lkReqRlseLoc_payload_txnAbt || (_zz_cntRlseReqWrLoc_0 < _zz_when_TxnManCS_l440_2)) || (_zz_cntRlseReqWrLoc_0 == 6'h0))) && (_zz_cntRlseReqLoc_0 < _zz_when_TxnManCS_l440)) || (_zz_lkReqRlseLoc_payload_txnTimeOut && (_zz_cntRlseReqLoc_0 < _zz_when_TxnManCS_l440_3)));
  assign lkReqRlseLoc_fire = (lkReqRlseLoc_valid && lkReqRlseLoc_ready);
  assign _zz_cntRlseReqLoc_0_1 = (_zz_cntRlseReqLoc_0 + 6'h01);
  assign lkReqRlseLoc_fire_1 = (lkReqRlseLoc_valid && lkReqRlseLoc_ready);
  assign when_TxnManCS_l456 = (lkReqRlseLoc_fire_1 && ((compLkRlseLoc_lkItem_lkType == LkT_wr) || (compLkRlseLoc_lkItem_lkType == LkT_raw)));
  assign _zz_cntRlseReqWrLoc_0_1 = (_zz_cntRlseReqWrLoc_0 + 6'h01);
  always @(*) begin
    compLkRlseRmt_stateNext = compLkRlseRmt_stateReg;
    case(compLkRlseRmt_stateReg)
      compLkRlseRmt_enumDef_CS_TXN : begin
        if(when_TxnManCS_l489) begin
          compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_RMT_LK_RLSE;
        end
      end
      compLkRlseRmt_enumDef_RMT_LK_RLSE : begin
        if(lkReqRlseRmt_fire) begin
          if(when_TxnManCS_l505) begin
            compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_RMT_WR;
          end else begin
            compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_CS_TXN;
          end
        end
      end
      compLkRlseRmt_enumDef_RMT_WR : begin
        if(io_wrRmt_fire) begin
          if(when_TxnManCS_l521) begin
            compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_CS_TXN;
          end
        end
      end
      default : begin
      end
    endcase
    if(compLkRlseRmt_wantStart) begin
      compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_CS_TXN;
    end
    if(compLkRlseRmt_wantKill) begin
      compLkRlseRmt_stateNext = compLkRlseRmt_enumDef_BOOT;
    end
  end

  assign _zz_when_TxnManCS_l489 = _zz__zz_when_TxnManCS_l489;
  assign when_TxnManCS_l489 = (((compLkRlseRmt_getAllLkResp && (_zz_lkReqRlseRmt_payload_txnAbt || _zz_when_TxnManCS_l489_1)) && (_zz_cntRlseReqRmt_0 < _zz_when_TxnManCS_l489)) || (_zz_lkReqRlseRmt_payload_txnTimeOut && (_zz_cntRlseReqRmt_0 < _zz_when_TxnManCS_l489_2)));
  assign lkReqRlseRmt_fire = (lkReqRlseRmt_valid && lkReqRlseRmt_ready);
  assign when_TxnManCS_l505 = (((compLkRlseRmt_lkItem_lkType == LkT_wr) || (compLkRlseRmt_lkItem_lkType == LkT_raw)) && (! _zz_lkReqRlseRmt_payload_txnAbt));
  assign _zz_350 = ({63'd0,1'b1} <<< compLkRlseRmt_curTxnId);
  assign _zz_cntRlseReqWrRmt_0 = (_zz__zz_cntRlseReqWrRmt_0 + 6'h01);
  assign _zz_cntRlseReqRmt_0_1 = (_zz_cntRlseReqRmt_0 + 6'h01);
  assign io_wrRmt_fire = (io_wrRmt_valid && io_wrRmt_ready);
  assign when_TxnManCS_l521 = (compLkRlseRmt_nBeat == _zz_when_TxnManCS_l521);
  assign _zz_cntRlseReqRmt_0_2 = (_zz_cntRlseReqRmt_0 + 6'h01);
  always @(*) begin
    compTimeOut_stateNext = compTimeOut_stateReg;
    case(compTimeOut_stateReg)
      compTimeOut_enumDef_IDLE : begin
        if(io_start) begin
          compTimeOut_stateNext = compTimeOut_enumDef_COUNT;
        end
      end
      compTimeOut_enumDef_COUNT : begin
        if(io_done) begin
          compTimeOut_stateNext = compTimeOut_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(compTimeOut_wantStart) begin
      compTimeOut_stateNext = compTimeOut_enumDef_IDLE;
    end
    if(compTimeOut_wantKill) begin
      compTimeOut_stateNext = compTimeOut_enumDef_BOOT;
    end
  end

  assign when_TxnManCS_l555 = (&cntTimeOut_0);
  assign when_TxnManCS_l555_1 = (&cntTimeOut_1);
  assign when_TxnManCS_l555_2 = (&cntTimeOut_2);
  assign when_TxnManCS_l555_3 = (&cntTimeOut_3);
  assign when_TxnManCS_l555_4 = (&cntTimeOut_4);
  assign when_TxnManCS_l555_5 = (&cntTimeOut_5);
  assign when_TxnManCS_l555_6 = (&cntTimeOut_6);
  assign when_TxnManCS_l555_7 = (&cntTimeOut_7);
  assign when_TxnManCS_l555_8 = (&cntTimeOut_8);
  assign when_TxnManCS_l555_9 = (&cntTimeOut_9);
  assign when_TxnManCS_l555_10 = (&cntTimeOut_10);
  assign when_TxnManCS_l555_11 = (&cntTimeOut_11);
  assign when_TxnManCS_l555_12 = (&cntTimeOut_12);
  assign when_TxnManCS_l555_13 = (&cntTimeOut_13);
  assign when_TxnManCS_l555_14 = (&cntTimeOut_14);
  assign when_TxnManCS_l555_15 = (&cntTimeOut_15);
  assign when_TxnManCS_l555_16 = (&cntTimeOut_16);
  assign when_TxnManCS_l555_17 = (&cntTimeOut_17);
  assign when_TxnManCS_l555_18 = (&cntTimeOut_18);
  assign when_TxnManCS_l555_19 = (&cntTimeOut_19);
  assign when_TxnManCS_l555_20 = (&cntTimeOut_20);
  assign when_TxnManCS_l555_21 = (&cntTimeOut_21);
  assign when_TxnManCS_l555_22 = (&cntTimeOut_22);
  assign when_TxnManCS_l555_23 = (&cntTimeOut_23);
  assign when_TxnManCS_l555_24 = (&cntTimeOut_24);
  assign when_TxnManCS_l555_25 = (&cntTimeOut_25);
  assign when_TxnManCS_l555_26 = (&cntTimeOut_26);
  assign when_TxnManCS_l555_27 = (&cntTimeOut_27);
  assign when_TxnManCS_l555_28 = (&cntTimeOut_28);
  assign when_TxnManCS_l555_29 = (&cntTimeOut_29);
  assign when_TxnManCS_l555_30 = (&cntTimeOut_30);
  assign when_TxnManCS_l555_31 = (&cntTimeOut_31);
  assign when_TxnManCS_l555_32 = (&cntTimeOut_32);
  assign when_TxnManCS_l555_33 = (&cntTimeOut_33);
  assign when_TxnManCS_l555_34 = (&cntTimeOut_34);
  assign when_TxnManCS_l555_35 = (&cntTimeOut_35);
  assign when_TxnManCS_l555_36 = (&cntTimeOut_36);
  assign when_TxnManCS_l555_37 = (&cntTimeOut_37);
  assign when_TxnManCS_l555_38 = (&cntTimeOut_38);
  assign when_TxnManCS_l555_39 = (&cntTimeOut_39);
  assign when_TxnManCS_l555_40 = (&cntTimeOut_40);
  assign when_TxnManCS_l555_41 = (&cntTimeOut_41);
  assign when_TxnManCS_l555_42 = (&cntTimeOut_42);
  assign when_TxnManCS_l555_43 = (&cntTimeOut_43);
  assign when_TxnManCS_l555_44 = (&cntTimeOut_44);
  assign when_TxnManCS_l555_45 = (&cntTimeOut_45);
  assign when_TxnManCS_l555_46 = (&cntTimeOut_46);
  assign when_TxnManCS_l555_47 = (&cntTimeOut_47);
  assign when_TxnManCS_l555_48 = (&cntTimeOut_48);
  assign when_TxnManCS_l555_49 = (&cntTimeOut_49);
  assign when_TxnManCS_l555_50 = (&cntTimeOut_50);
  assign when_TxnManCS_l555_51 = (&cntTimeOut_51);
  assign when_TxnManCS_l555_52 = (&cntTimeOut_52);
  assign when_TxnManCS_l555_53 = (&cntTimeOut_53);
  assign when_TxnManCS_l555_54 = (&cntTimeOut_54);
  assign when_TxnManCS_l555_55 = (&cntTimeOut_55);
  assign when_TxnManCS_l555_56 = (&cntTimeOut_56);
  assign when_TxnManCS_l555_57 = (&cntTimeOut_57);
  assign when_TxnManCS_l555_58 = (&cntTimeOut_58);
  assign when_TxnManCS_l555_59 = (&cntTimeOut_59);
  assign when_TxnManCS_l555_60 = (&cntTimeOut_60);
  assign when_TxnManCS_l555_61 = (&cntTimeOut_61);
  assign when_TxnManCS_l555_62 = (&cntTimeOut_62);
  assign when_TxnManCS_l555_63 = (&cntTimeOut_63);
  always @(*) begin
    compLoadTxn_stateNext = compLoadTxn_stateReg;
    case(compLoadTxn_stateReg)
      compLoadTxn_enumDef_IDLE : begin
        if(io_start) begin
          compLoadTxn_stateNext = compLoadTxn_enumDef_CS_TXN;
        end
      end
      compLoadTxn_enumDef_CS_TXN : begin
        if(when_TxnManCS_l621) begin
          compLoadTxn_stateNext = compLoadTxn_enumDef_RD_CMDAXI;
        end
      end
      compLoadTxn_enumDef_RD_CMDAXI : begin
        if(io_cmdAxi_ar_fire) begin
          compLoadTxn_stateNext = compLoadTxn_enumDef_LD_TXN;
        end
      end
      compLoadTxn_enumDef_LD_TXN : begin
        if(compLoadTxn_cntTxnWord_willOverflow) begin
          if(when_TxnManCS_l665) begin
            compLoadTxn_stateNext = compLoadTxn_enumDef_IDLE;
          end else begin
            compLoadTxn_stateNext = compLoadTxn_enumDef_CS_TXN;
          end
        end
      end
      default : begin
      end
    endcase
    if(compLoadTxn_wantStart) begin
      compLoadTxn_stateNext = compLoadTxn_enumDef_IDLE;
    end
    if(compLoadTxn_wantKill) begin
      compLoadTxn_stateNext = compLoadTxn_enumDef_BOOT;
    end
  end

  assign when_TxnManCS_l621 = _zz_when_TxnManCS_l621;
  assign _zz_351 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign io_cmdAxi_ar_fire = (io_cmdAxi_ar_valid && io_cmdAxi_ar_ready);
  assign io_cmdAxi_r_fire_2 = (io_cmdAxi_r_valid && io_cmdAxi_r_ready);
  assign _zz_353 = compLoadTxn_txnBuff[27 : 26];
  assign _zz_352 = _zz_353;
  assign _zz_354 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_355 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_356 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_357 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_358 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_359 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_360 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_361 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_362 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_363 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_364 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_365 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_366 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_367 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_368 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_369 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_370 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_371 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_372 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_373 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_374 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_375 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_376 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_377 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_378 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign _zz_379 = ({63'd0,1'b1} <<< compLoadTxn_curTxnId);
  assign when_TxnManCS_l665 = (compLoadTxn_cntTxn == _zz_when_TxnManCS_l665);
  always @(*) begin
    clkCnt_stateNext = clkCnt_stateReg;
    case(clkCnt_stateReg)
      clkCnt_enumDef_IDLE : begin
        if(io_start) begin
          clkCnt_stateNext = clkCnt_enumDef_CNT;
        end
      end
      clkCnt_enumDef_CNT : begin
        if(io_done) begin
          clkCnt_stateNext = clkCnt_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(clkCnt_wantStart) begin
      clkCnt_stateNext = clkCnt_enumDef_IDLE;
    end
    if(clkCnt_wantKill) begin
      clkCnt_stateNext = clkCnt_enumDef_BOOT;
    end
  end

  always @(posedge clk) begin
    if(!resetn) begin
      io_done <= 1'b0;
      io_cntTxnCmt <= 32'h0;
      io_cntTxnAbt <= 32'h0;
      io_cntTxnLd <= 32'h0;
      io_cntLockLoc <= 32'h0;
      io_cntLockRmt <= 32'h0;
      io_cntLockDenyLoc <= 32'h0;
      io_cntLockDenyRmt <= 32'h0;
      io_cntClk <= 32'h0;
      streamArbiter_8_io_output_rValid <= 1'b0;
      streamArbiter_8_io_output_s2mPipe_rValid <= 1'b0;
      streamArbiter_9_io_output_rValid <= 1'b0;
      streamArbiter_9_io_output_s2mPipe_rValid <= 1'b0;
      cntLkReqLoc_0 <= 6'h0;
      cntLkReqLoc_1 <= 6'h0;
      cntLkReqLoc_2 <= 6'h0;
      cntLkReqLoc_3 <= 6'h0;
      cntLkReqLoc_4 <= 6'h0;
      cntLkReqLoc_5 <= 6'h0;
      cntLkReqLoc_6 <= 6'h0;
      cntLkReqLoc_7 <= 6'h0;
      cntLkReqLoc_8 <= 6'h0;
      cntLkReqLoc_9 <= 6'h0;
      cntLkReqLoc_10 <= 6'h0;
      cntLkReqLoc_11 <= 6'h0;
      cntLkReqLoc_12 <= 6'h0;
      cntLkReqLoc_13 <= 6'h0;
      cntLkReqLoc_14 <= 6'h0;
      cntLkReqLoc_15 <= 6'h0;
      cntLkReqLoc_16 <= 6'h0;
      cntLkReqLoc_17 <= 6'h0;
      cntLkReqLoc_18 <= 6'h0;
      cntLkReqLoc_19 <= 6'h0;
      cntLkReqLoc_20 <= 6'h0;
      cntLkReqLoc_21 <= 6'h0;
      cntLkReqLoc_22 <= 6'h0;
      cntLkReqLoc_23 <= 6'h0;
      cntLkReqLoc_24 <= 6'h0;
      cntLkReqLoc_25 <= 6'h0;
      cntLkReqLoc_26 <= 6'h0;
      cntLkReqLoc_27 <= 6'h0;
      cntLkReqLoc_28 <= 6'h0;
      cntLkReqLoc_29 <= 6'h0;
      cntLkReqLoc_30 <= 6'h0;
      cntLkReqLoc_31 <= 6'h0;
      cntLkReqLoc_32 <= 6'h0;
      cntLkReqLoc_33 <= 6'h0;
      cntLkReqLoc_34 <= 6'h0;
      cntLkReqLoc_35 <= 6'h0;
      cntLkReqLoc_36 <= 6'h0;
      cntLkReqLoc_37 <= 6'h0;
      cntLkReqLoc_38 <= 6'h0;
      cntLkReqLoc_39 <= 6'h0;
      cntLkReqLoc_40 <= 6'h0;
      cntLkReqLoc_41 <= 6'h0;
      cntLkReqLoc_42 <= 6'h0;
      cntLkReqLoc_43 <= 6'h0;
      cntLkReqLoc_44 <= 6'h0;
      cntLkReqLoc_45 <= 6'h0;
      cntLkReqLoc_46 <= 6'h0;
      cntLkReqLoc_47 <= 6'h0;
      cntLkReqLoc_48 <= 6'h0;
      cntLkReqLoc_49 <= 6'h0;
      cntLkReqLoc_50 <= 6'h0;
      cntLkReqLoc_51 <= 6'h0;
      cntLkReqLoc_52 <= 6'h0;
      cntLkReqLoc_53 <= 6'h0;
      cntLkReqLoc_54 <= 6'h0;
      cntLkReqLoc_55 <= 6'h0;
      cntLkReqLoc_56 <= 6'h0;
      cntLkReqLoc_57 <= 6'h0;
      cntLkReqLoc_58 <= 6'h0;
      cntLkReqLoc_59 <= 6'h0;
      cntLkReqLoc_60 <= 6'h0;
      cntLkReqLoc_61 <= 6'h0;
      cntLkReqLoc_62 <= 6'h0;
      cntLkReqLoc_63 <= 6'h0;
      cntLkReqRmt_0 <= 6'h0;
      cntLkReqRmt_1 <= 6'h0;
      cntLkReqRmt_2 <= 6'h0;
      cntLkReqRmt_3 <= 6'h0;
      cntLkReqRmt_4 <= 6'h0;
      cntLkReqRmt_5 <= 6'h0;
      cntLkReqRmt_6 <= 6'h0;
      cntLkReqRmt_7 <= 6'h0;
      cntLkReqRmt_8 <= 6'h0;
      cntLkReqRmt_9 <= 6'h0;
      cntLkReqRmt_10 <= 6'h0;
      cntLkReqRmt_11 <= 6'h0;
      cntLkReqRmt_12 <= 6'h0;
      cntLkReqRmt_13 <= 6'h0;
      cntLkReqRmt_14 <= 6'h0;
      cntLkReqRmt_15 <= 6'h0;
      cntLkReqRmt_16 <= 6'h0;
      cntLkReqRmt_17 <= 6'h0;
      cntLkReqRmt_18 <= 6'h0;
      cntLkReqRmt_19 <= 6'h0;
      cntLkReqRmt_20 <= 6'h0;
      cntLkReqRmt_21 <= 6'h0;
      cntLkReqRmt_22 <= 6'h0;
      cntLkReqRmt_23 <= 6'h0;
      cntLkReqRmt_24 <= 6'h0;
      cntLkReqRmt_25 <= 6'h0;
      cntLkReqRmt_26 <= 6'h0;
      cntLkReqRmt_27 <= 6'h0;
      cntLkReqRmt_28 <= 6'h0;
      cntLkReqRmt_29 <= 6'h0;
      cntLkReqRmt_30 <= 6'h0;
      cntLkReqRmt_31 <= 6'h0;
      cntLkReqRmt_32 <= 6'h0;
      cntLkReqRmt_33 <= 6'h0;
      cntLkReqRmt_34 <= 6'h0;
      cntLkReqRmt_35 <= 6'h0;
      cntLkReqRmt_36 <= 6'h0;
      cntLkReqRmt_37 <= 6'h0;
      cntLkReqRmt_38 <= 6'h0;
      cntLkReqRmt_39 <= 6'h0;
      cntLkReqRmt_40 <= 6'h0;
      cntLkReqRmt_41 <= 6'h0;
      cntLkReqRmt_42 <= 6'h0;
      cntLkReqRmt_43 <= 6'h0;
      cntLkReqRmt_44 <= 6'h0;
      cntLkReqRmt_45 <= 6'h0;
      cntLkReqRmt_46 <= 6'h0;
      cntLkReqRmt_47 <= 6'h0;
      cntLkReqRmt_48 <= 6'h0;
      cntLkReqRmt_49 <= 6'h0;
      cntLkReqRmt_50 <= 6'h0;
      cntLkReqRmt_51 <= 6'h0;
      cntLkReqRmt_52 <= 6'h0;
      cntLkReqRmt_53 <= 6'h0;
      cntLkReqRmt_54 <= 6'h0;
      cntLkReqRmt_55 <= 6'h0;
      cntLkReqRmt_56 <= 6'h0;
      cntLkReqRmt_57 <= 6'h0;
      cntLkReqRmt_58 <= 6'h0;
      cntLkReqRmt_59 <= 6'h0;
      cntLkReqRmt_60 <= 6'h0;
      cntLkReqRmt_61 <= 6'h0;
      cntLkReqRmt_62 <= 6'h0;
      cntLkReqRmt_63 <= 6'h0;
      cntLkRespLoc_0 <= 6'h0;
      cntLkRespLoc_1 <= 6'h0;
      cntLkRespLoc_2 <= 6'h0;
      cntLkRespLoc_3 <= 6'h0;
      cntLkRespLoc_4 <= 6'h0;
      cntLkRespLoc_5 <= 6'h0;
      cntLkRespLoc_6 <= 6'h0;
      cntLkRespLoc_7 <= 6'h0;
      cntLkRespLoc_8 <= 6'h0;
      cntLkRespLoc_9 <= 6'h0;
      cntLkRespLoc_10 <= 6'h0;
      cntLkRespLoc_11 <= 6'h0;
      cntLkRespLoc_12 <= 6'h0;
      cntLkRespLoc_13 <= 6'h0;
      cntLkRespLoc_14 <= 6'h0;
      cntLkRespLoc_15 <= 6'h0;
      cntLkRespLoc_16 <= 6'h0;
      cntLkRespLoc_17 <= 6'h0;
      cntLkRespLoc_18 <= 6'h0;
      cntLkRespLoc_19 <= 6'h0;
      cntLkRespLoc_20 <= 6'h0;
      cntLkRespLoc_21 <= 6'h0;
      cntLkRespLoc_22 <= 6'h0;
      cntLkRespLoc_23 <= 6'h0;
      cntLkRespLoc_24 <= 6'h0;
      cntLkRespLoc_25 <= 6'h0;
      cntLkRespLoc_26 <= 6'h0;
      cntLkRespLoc_27 <= 6'h0;
      cntLkRespLoc_28 <= 6'h0;
      cntLkRespLoc_29 <= 6'h0;
      cntLkRespLoc_30 <= 6'h0;
      cntLkRespLoc_31 <= 6'h0;
      cntLkRespLoc_32 <= 6'h0;
      cntLkRespLoc_33 <= 6'h0;
      cntLkRespLoc_34 <= 6'h0;
      cntLkRespLoc_35 <= 6'h0;
      cntLkRespLoc_36 <= 6'h0;
      cntLkRespLoc_37 <= 6'h0;
      cntLkRespLoc_38 <= 6'h0;
      cntLkRespLoc_39 <= 6'h0;
      cntLkRespLoc_40 <= 6'h0;
      cntLkRespLoc_41 <= 6'h0;
      cntLkRespLoc_42 <= 6'h0;
      cntLkRespLoc_43 <= 6'h0;
      cntLkRespLoc_44 <= 6'h0;
      cntLkRespLoc_45 <= 6'h0;
      cntLkRespLoc_46 <= 6'h0;
      cntLkRespLoc_47 <= 6'h0;
      cntLkRespLoc_48 <= 6'h0;
      cntLkRespLoc_49 <= 6'h0;
      cntLkRespLoc_50 <= 6'h0;
      cntLkRespLoc_51 <= 6'h0;
      cntLkRespLoc_52 <= 6'h0;
      cntLkRespLoc_53 <= 6'h0;
      cntLkRespLoc_54 <= 6'h0;
      cntLkRespLoc_55 <= 6'h0;
      cntLkRespLoc_56 <= 6'h0;
      cntLkRespLoc_57 <= 6'h0;
      cntLkRespLoc_58 <= 6'h0;
      cntLkRespLoc_59 <= 6'h0;
      cntLkRespLoc_60 <= 6'h0;
      cntLkRespLoc_61 <= 6'h0;
      cntLkRespLoc_62 <= 6'h0;
      cntLkRespLoc_63 <= 6'h0;
      cntLkRespRmt_0 <= 6'h0;
      cntLkRespRmt_1 <= 6'h0;
      cntLkRespRmt_2 <= 6'h0;
      cntLkRespRmt_3 <= 6'h0;
      cntLkRespRmt_4 <= 6'h0;
      cntLkRespRmt_5 <= 6'h0;
      cntLkRespRmt_6 <= 6'h0;
      cntLkRespRmt_7 <= 6'h0;
      cntLkRespRmt_8 <= 6'h0;
      cntLkRespRmt_9 <= 6'h0;
      cntLkRespRmt_10 <= 6'h0;
      cntLkRespRmt_11 <= 6'h0;
      cntLkRespRmt_12 <= 6'h0;
      cntLkRespRmt_13 <= 6'h0;
      cntLkRespRmt_14 <= 6'h0;
      cntLkRespRmt_15 <= 6'h0;
      cntLkRespRmt_16 <= 6'h0;
      cntLkRespRmt_17 <= 6'h0;
      cntLkRespRmt_18 <= 6'h0;
      cntLkRespRmt_19 <= 6'h0;
      cntLkRespRmt_20 <= 6'h0;
      cntLkRespRmt_21 <= 6'h0;
      cntLkRespRmt_22 <= 6'h0;
      cntLkRespRmt_23 <= 6'h0;
      cntLkRespRmt_24 <= 6'h0;
      cntLkRespRmt_25 <= 6'h0;
      cntLkRespRmt_26 <= 6'h0;
      cntLkRespRmt_27 <= 6'h0;
      cntLkRespRmt_28 <= 6'h0;
      cntLkRespRmt_29 <= 6'h0;
      cntLkRespRmt_30 <= 6'h0;
      cntLkRespRmt_31 <= 6'h0;
      cntLkRespRmt_32 <= 6'h0;
      cntLkRespRmt_33 <= 6'h0;
      cntLkRespRmt_34 <= 6'h0;
      cntLkRespRmt_35 <= 6'h0;
      cntLkRespRmt_36 <= 6'h0;
      cntLkRespRmt_37 <= 6'h0;
      cntLkRespRmt_38 <= 6'h0;
      cntLkRespRmt_39 <= 6'h0;
      cntLkRespRmt_40 <= 6'h0;
      cntLkRespRmt_41 <= 6'h0;
      cntLkRespRmt_42 <= 6'h0;
      cntLkRespRmt_43 <= 6'h0;
      cntLkRespRmt_44 <= 6'h0;
      cntLkRespRmt_45 <= 6'h0;
      cntLkRespRmt_46 <= 6'h0;
      cntLkRespRmt_47 <= 6'h0;
      cntLkRespRmt_48 <= 6'h0;
      cntLkRespRmt_49 <= 6'h0;
      cntLkRespRmt_50 <= 6'h0;
      cntLkRespRmt_51 <= 6'h0;
      cntLkRespRmt_52 <= 6'h0;
      cntLkRespRmt_53 <= 6'h0;
      cntLkRespRmt_54 <= 6'h0;
      cntLkRespRmt_55 <= 6'h0;
      cntLkRespRmt_56 <= 6'h0;
      cntLkRespRmt_57 <= 6'h0;
      cntLkRespRmt_58 <= 6'h0;
      cntLkRespRmt_59 <= 6'h0;
      cntLkRespRmt_60 <= 6'h0;
      cntLkRespRmt_61 <= 6'h0;
      cntLkRespRmt_62 <= 6'h0;
      cntLkRespRmt_63 <= 6'h0;
      cntLkHoldLoc_0 <= 6'h0;
      cntLkHoldLoc_1 <= 6'h0;
      cntLkHoldLoc_2 <= 6'h0;
      cntLkHoldLoc_3 <= 6'h0;
      cntLkHoldLoc_4 <= 6'h0;
      cntLkHoldLoc_5 <= 6'h0;
      cntLkHoldLoc_6 <= 6'h0;
      cntLkHoldLoc_7 <= 6'h0;
      cntLkHoldLoc_8 <= 6'h0;
      cntLkHoldLoc_9 <= 6'h0;
      cntLkHoldLoc_10 <= 6'h0;
      cntLkHoldLoc_11 <= 6'h0;
      cntLkHoldLoc_12 <= 6'h0;
      cntLkHoldLoc_13 <= 6'h0;
      cntLkHoldLoc_14 <= 6'h0;
      cntLkHoldLoc_15 <= 6'h0;
      cntLkHoldLoc_16 <= 6'h0;
      cntLkHoldLoc_17 <= 6'h0;
      cntLkHoldLoc_18 <= 6'h0;
      cntLkHoldLoc_19 <= 6'h0;
      cntLkHoldLoc_20 <= 6'h0;
      cntLkHoldLoc_21 <= 6'h0;
      cntLkHoldLoc_22 <= 6'h0;
      cntLkHoldLoc_23 <= 6'h0;
      cntLkHoldLoc_24 <= 6'h0;
      cntLkHoldLoc_25 <= 6'h0;
      cntLkHoldLoc_26 <= 6'h0;
      cntLkHoldLoc_27 <= 6'h0;
      cntLkHoldLoc_28 <= 6'h0;
      cntLkHoldLoc_29 <= 6'h0;
      cntLkHoldLoc_30 <= 6'h0;
      cntLkHoldLoc_31 <= 6'h0;
      cntLkHoldLoc_32 <= 6'h0;
      cntLkHoldLoc_33 <= 6'h0;
      cntLkHoldLoc_34 <= 6'h0;
      cntLkHoldLoc_35 <= 6'h0;
      cntLkHoldLoc_36 <= 6'h0;
      cntLkHoldLoc_37 <= 6'h0;
      cntLkHoldLoc_38 <= 6'h0;
      cntLkHoldLoc_39 <= 6'h0;
      cntLkHoldLoc_40 <= 6'h0;
      cntLkHoldLoc_41 <= 6'h0;
      cntLkHoldLoc_42 <= 6'h0;
      cntLkHoldLoc_43 <= 6'h0;
      cntLkHoldLoc_44 <= 6'h0;
      cntLkHoldLoc_45 <= 6'h0;
      cntLkHoldLoc_46 <= 6'h0;
      cntLkHoldLoc_47 <= 6'h0;
      cntLkHoldLoc_48 <= 6'h0;
      cntLkHoldLoc_49 <= 6'h0;
      cntLkHoldLoc_50 <= 6'h0;
      cntLkHoldLoc_51 <= 6'h0;
      cntLkHoldLoc_52 <= 6'h0;
      cntLkHoldLoc_53 <= 6'h0;
      cntLkHoldLoc_54 <= 6'h0;
      cntLkHoldLoc_55 <= 6'h0;
      cntLkHoldLoc_56 <= 6'h0;
      cntLkHoldLoc_57 <= 6'h0;
      cntLkHoldLoc_58 <= 6'h0;
      cntLkHoldLoc_59 <= 6'h0;
      cntLkHoldLoc_60 <= 6'h0;
      cntLkHoldLoc_61 <= 6'h0;
      cntLkHoldLoc_62 <= 6'h0;
      cntLkHoldLoc_63 <= 6'h0;
      cntLkHoldRmt_0 <= 6'h0;
      cntLkHoldRmt_1 <= 6'h0;
      cntLkHoldRmt_2 <= 6'h0;
      cntLkHoldRmt_3 <= 6'h0;
      cntLkHoldRmt_4 <= 6'h0;
      cntLkHoldRmt_5 <= 6'h0;
      cntLkHoldRmt_6 <= 6'h0;
      cntLkHoldRmt_7 <= 6'h0;
      cntLkHoldRmt_8 <= 6'h0;
      cntLkHoldRmt_9 <= 6'h0;
      cntLkHoldRmt_10 <= 6'h0;
      cntLkHoldRmt_11 <= 6'h0;
      cntLkHoldRmt_12 <= 6'h0;
      cntLkHoldRmt_13 <= 6'h0;
      cntLkHoldRmt_14 <= 6'h0;
      cntLkHoldRmt_15 <= 6'h0;
      cntLkHoldRmt_16 <= 6'h0;
      cntLkHoldRmt_17 <= 6'h0;
      cntLkHoldRmt_18 <= 6'h0;
      cntLkHoldRmt_19 <= 6'h0;
      cntLkHoldRmt_20 <= 6'h0;
      cntLkHoldRmt_21 <= 6'h0;
      cntLkHoldRmt_22 <= 6'h0;
      cntLkHoldRmt_23 <= 6'h0;
      cntLkHoldRmt_24 <= 6'h0;
      cntLkHoldRmt_25 <= 6'h0;
      cntLkHoldRmt_26 <= 6'h0;
      cntLkHoldRmt_27 <= 6'h0;
      cntLkHoldRmt_28 <= 6'h0;
      cntLkHoldRmt_29 <= 6'h0;
      cntLkHoldRmt_30 <= 6'h0;
      cntLkHoldRmt_31 <= 6'h0;
      cntLkHoldRmt_32 <= 6'h0;
      cntLkHoldRmt_33 <= 6'h0;
      cntLkHoldRmt_34 <= 6'h0;
      cntLkHoldRmt_35 <= 6'h0;
      cntLkHoldRmt_36 <= 6'h0;
      cntLkHoldRmt_37 <= 6'h0;
      cntLkHoldRmt_38 <= 6'h0;
      cntLkHoldRmt_39 <= 6'h0;
      cntLkHoldRmt_40 <= 6'h0;
      cntLkHoldRmt_41 <= 6'h0;
      cntLkHoldRmt_42 <= 6'h0;
      cntLkHoldRmt_43 <= 6'h0;
      cntLkHoldRmt_44 <= 6'h0;
      cntLkHoldRmt_45 <= 6'h0;
      cntLkHoldRmt_46 <= 6'h0;
      cntLkHoldRmt_47 <= 6'h0;
      cntLkHoldRmt_48 <= 6'h0;
      cntLkHoldRmt_49 <= 6'h0;
      cntLkHoldRmt_50 <= 6'h0;
      cntLkHoldRmt_51 <= 6'h0;
      cntLkHoldRmt_52 <= 6'h0;
      cntLkHoldRmt_53 <= 6'h0;
      cntLkHoldRmt_54 <= 6'h0;
      cntLkHoldRmt_55 <= 6'h0;
      cntLkHoldRmt_56 <= 6'h0;
      cntLkHoldRmt_57 <= 6'h0;
      cntLkHoldRmt_58 <= 6'h0;
      cntLkHoldRmt_59 <= 6'h0;
      cntLkHoldRmt_60 <= 6'h0;
      cntLkHoldRmt_61 <= 6'h0;
      cntLkHoldRmt_62 <= 6'h0;
      cntLkHoldRmt_63 <= 6'h0;
      cntLkWaitLoc_0 <= 6'h0;
      cntLkWaitLoc_1 <= 6'h0;
      cntLkWaitLoc_2 <= 6'h0;
      cntLkWaitLoc_3 <= 6'h0;
      cntLkWaitLoc_4 <= 6'h0;
      cntLkWaitLoc_5 <= 6'h0;
      cntLkWaitLoc_6 <= 6'h0;
      cntLkWaitLoc_7 <= 6'h0;
      cntLkWaitLoc_8 <= 6'h0;
      cntLkWaitLoc_9 <= 6'h0;
      cntLkWaitLoc_10 <= 6'h0;
      cntLkWaitLoc_11 <= 6'h0;
      cntLkWaitLoc_12 <= 6'h0;
      cntLkWaitLoc_13 <= 6'h0;
      cntLkWaitLoc_14 <= 6'h0;
      cntLkWaitLoc_15 <= 6'h0;
      cntLkWaitLoc_16 <= 6'h0;
      cntLkWaitLoc_17 <= 6'h0;
      cntLkWaitLoc_18 <= 6'h0;
      cntLkWaitLoc_19 <= 6'h0;
      cntLkWaitLoc_20 <= 6'h0;
      cntLkWaitLoc_21 <= 6'h0;
      cntLkWaitLoc_22 <= 6'h0;
      cntLkWaitLoc_23 <= 6'h0;
      cntLkWaitLoc_24 <= 6'h0;
      cntLkWaitLoc_25 <= 6'h0;
      cntLkWaitLoc_26 <= 6'h0;
      cntLkWaitLoc_27 <= 6'h0;
      cntLkWaitLoc_28 <= 6'h0;
      cntLkWaitLoc_29 <= 6'h0;
      cntLkWaitLoc_30 <= 6'h0;
      cntLkWaitLoc_31 <= 6'h0;
      cntLkWaitLoc_32 <= 6'h0;
      cntLkWaitLoc_33 <= 6'h0;
      cntLkWaitLoc_34 <= 6'h0;
      cntLkWaitLoc_35 <= 6'h0;
      cntLkWaitLoc_36 <= 6'h0;
      cntLkWaitLoc_37 <= 6'h0;
      cntLkWaitLoc_38 <= 6'h0;
      cntLkWaitLoc_39 <= 6'h0;
      cntLkWaitLoc_40 <= 6'h0;
      cntLkWaitLoc_41 <= 6'h0;
      cntLkWaitLoc_42 <= 6'h0;
      cntLkWaitLoc_43 <= 6'h0;
      cntLkWaitLoc_44 <= 6'h0;
      cntLkWaitLoc_45 <= 6'h0;
      cntLkWaitLoc_46 <= 6'h0;
      cntLkWaitLoc_47 <= 6'h0;
      cntLkWaitLoc_48 <= 6'h0;
      cntLkWaitLoc_49 <= 6'h0;
      cntLkWaitLoc_50 <= 6'h0;
      cntLkWaitLoc_51 <= 6'h0;
      cntLkWaitLoc_52 <= 6'h0;
      cntLkWaitLoc_53 <= 6'h0;
      cntLkWaitLoc_54 <= 6'h0;
      cntLkWaitLoc_55 <= 6'h0;
      cntLkWaitLoc_56 <= 6'h0;
      cntLkWaitLoc_57 <= 6'h0;
      cntLkWaitLoc_58 <= 6'h0;
      cntLkWaitLoc_59 <= 6'h0;
      cntLkWaitLoc_60 <= 6'h0;
      cntLkWaitLoc_61 <= 6'h0;
      cntLkWaitLoc_62 <= 6'h0;
      cntLkWaitLoc_63 <= 6'h0;
      cntLkWaitRmt_0 <= 6'h0;
      cntLkWaitRmt_1 <= 6'h0;
      cntLkWaitRmt_2 <= 6'h0;
      cntLkWaitRmt_3 <= 6'h0;
      cntLkWaitRmt_4 <= 6'h0;
      cntLkWaitRmt_5 <= 6'h0;
      cntLkWaitRmt_6 <= 6'h0;
      cntLkWaitRmt_7 <= 6'h0;
      cntLkWaitRmt_8 <= 6'h0;
      cntLkWaitRmt_9 <= 6'h0;
      cntLkWaitRmt_10 <= 6'h0;
      cntLkWaitRmt_11 <= 6'h0;
      cntLkWaitRmt_12 <= 6'h0;
      cntLkWaitRmt_13 <= 6'h0;
      cntLkWaitRmt_14 <= 6'h0;
      cntLkWaitRmt_15 <= 6'h0;
      cntLkWaitRmt_16 <= 6'h0;
      cntLkWaitRmt_17 <= 6'h0;
      cntLkWaitRmt_18 <= 6'h0;
      cntLkWaitRmt_19 <= 6'h0;
      cntLkWaitRmt_20 <= 6'h0;
      cntLkWaitRmt_21 <= 6'h0;
      cntLkWaitRmt_22 <= 6'h0;
      cntLkWaitRmt_23 <= 6'h0;
      cntLkWaitRmt_24 <= 6'h0;
      cntLkWaitRmt_25 <= 6'h0;
      cntLkWaitRmt_26 <= 6'h0;
      cntLkWaitRmt_27 <= 6'h0;
      cntLkWaitRmt_28 <= 6'h0;
      cntLkWaitRmt_29 <= 6'h0;
      cntLkWaitRmt_30 <= 6'h0;
      cntLkWaitRmt_31 <= 6'h0;
      cntLkWaitRmt_32 <= 6'h0;
      cntLkWaitRmt_33 <= 6'h0;
      cntLkWaitRmt_34 <= 6'h0;
      cntLkWaitRmt_35 <= 6'h0;
      cntLkWaitRmt_36 <= 6'h0;
      cntLkWaitRmt_37 <= 6'h0;
      cntLkWaitRmt_38 <= 6'h0;
      cntLkWaitRmt_39 <= 6'h0;
      cntLkWaitRmt_40 <= 6'h0;
      cntLkWaitRmt_41 <= 6'h0;
      cntLkWaitRmt_42 <= 6'h0;
      cntLkWaitRmt_43 <= 6'h0;
      cntLkWaitRmt_44 <= 6'h0;
      cntLkWaitRmt_45 <= 6'h0;
      cntLkWaitRmt_46 <= 6'h0;
      cntLkWaitRmt_47 <= 6'h0;
      cntLkWaitRmt_48 <= 6'h0;
      cntLkWaitRmt_49 <= 6'h0;
      cntLkWaitRmt_50 <= 6'h0;
      cntLkWaitRmt_51 <= 6'h0;
      cntLkWaitRmt_52 <= 6'h0;
      cntLkWaitRmt_53 <= 6'h0;
      cntLkWaitRmt_54 <= 6'h0;
      cntLkWaitRmt_55 <= 6'h0;
      cntLkWaitRmt_56 <= 6'h0;
      cntLkWaitRmt_57 <= 6'h0;
      cntLkWaitRmt_58 <= 6'h0;
      cntLkWaitRmt_59 <= 6'h0;
      cntLkWaitRmt_60 <= 6'h0;
      cntLkWaitRmt_61 <= 6'h0;
      cntLkWaitRmt_62 <= 6'h0;
      cntLkWaitRmt_63 <= 6'h0;
      cntLkReqWrLoc_0 <= 6'h0;
      cntLkReqWrLoc_1 <= 6'h0;
      cntLkReqWrLoc_2 <= 6'h0;
      cntLkReqWrLoc_3 <= 6'h0;
      cntLkReqWrLoc_4 <= 6'h0;
      cntLkReqWrLoc_5 <= 6'h0;
      cntLkReqWrLoc_6 <= 6'h0;
      cntLkReqWrLoc_7 <= 6'h0;
      cntLkReqWrLoc_8 <= 6'h0;
      cntLkReqWrLoc_9 <= 6'h0;
      cntLkReqWrLoc_10 <= 6'h0;
      cntLkReqWrLoc_11 <= 6'h0;
      cntLkReqWrLoc_12 <= 6'h0;
      cntLkReqWrLoc_13 <= 6'h0;
      cntLkReqWrLoc_14 <= 6'h0;
      cntLkReqWrLoc_15 <= 6'h0;
      cntLkReqWrLoc_16 <= 6'h0;
      cntLkReqWrLoc_17 <= 6'h0;
      cntLkReqWrLoc_18 <= 6'h0;
      cntLkReqWrLoc_19 <= 6'h0;
      cntLkReqWrLoc_20 <= 6'h0;
      cntLkReqWrLoc_21 <= 6'h0;
      cntLkReqWrLoc_22 <= 6'h0;
      cntLkReqWrLoc_23 <= 6'h0;
      cntLkReqWrLoc_24 <= 6'h0;
      cntLkReqWrLoc_25 <= 6'h0;
      cntLkReqWrLoc_26 <= 6'h0;
      cntLkReqWrLoc_27 <= 6'h0;
      cntLkReqWrLoc_28 <= 6'h0;
      cntLkReqWrLoc_29 <= 6'h0;
      cntLkReqWrLoc_30 <= 6'h0;
      cntLkReqWrLoc_31 <= 6'h0;
      cntLkReqWrLoc_32 <= 6'h0;
      cntLkReqWrLoc_33 <= 6'h0;
      cntLkReqWrLoc_34 <= 6'h0;
      cntLkReqWrLoc_35 <= 6'h0;
      cntLkReqWrLoc_36 <= 6'h0;
      cntLkReqWrLoc_37 <= 6'h0;
      cntLkReqWrLoc_38 <= 6'h0;
      cntLkReqWrLoc_39 <= 6'h0;
      cntLkReqWrLoc_40 <= 6'h0;
      cntLkReqWrLoc_41 <= 6'h0;
      cntLkReqWrLoc_42 <= 6'h0;
      cntLkReqWrLoc_43 <= 6'h0;
      cntLkReqWrLoc_44 <= 6'h0;
      cntLkReqWrLoc_45 <= 6'h0;
      cntLkReqWrLoc_46 <= 6'h0;
      cntLkReqWrLoc_47 <= 6'h0;
      cntLkReqWrLoc_48 <= 6'h0;
      cntLkReqWrLoc_49 <= 6'h0;
      cntLkReqWrLoc_50 <= 6'h0;
      cntLkReqWrLoc_51 <= 6'h0;
      cntLkReqWrLoc_52 <= 6'h0;
      cntLkReqWrLoc_53 <= 6'h0;
      cntLkReqWrLoc_54 <= 6'h0;
      cntLkReqWrLoc_55 <= 6'h0;
      cntLkReqWrLoc_56 <= 6'h0;
      cntLkReqWrLoc_57 <= 6'h0;
      cntLkReqWrLoc_58 <= 6'h0;
      cntLkReqWrLoc_59 <= 6'h0;
      cntLkReqWrLoc_60 <= 6'h0;
      cntLkReqWrLoc_61 <= 6'h0;
      cntLkReqWrLoc_62 <= 6'h0;
      cntLkReqWrLoc_63 <= 6'h0;
      cntLkReqWrRmt_0 <= 6'h0;
      cntLkReqWrRmt_1 <= 6'h0;
      cntLkReqWrRmt_2 <= 6'h0;
      cntLkReqWrRmt_3 <= 6'h0;
      cntLkReqWrRmt_4 <= 6'h0;
      cntLkReqWrRmt_5 <= 6'h0;
      cntLkReqWrRmt_6 <= 6'h0;
      cntLkReqWrRmt_7 <= 6'h0;
      cntLkReqWrRmt_8 <= 6'h0;
      cntLkReqWrRmt_9 <= 6'h0;
      cntLkReqWrRmt_10 <= 6'h0;
      cntLkReqWrRmt_11 <= 6'h0;
      cntLkReqWrRmt_12 <= 6'h0;
      cntLkReqWrRmt_13 <= 6'h0;
      cntLkReqWrRmt_14 <= 6'h0;
      cntLkReqWrRmt_15 <= 6'h0;
      cntLkReqWrRmt_16 <= 6'h0;
      cntLkReqWrRmt_17 <= 6'h0;
      cntLkReqWrRmt_18 <= 6'h0;
      cntLkReqWrRmt_19 <= 6'h0;
      cntLkReqWrRmt_20 <= 6'h0;
      cntLkReqWrRmt_21 <= 6'h0;
      cntLkReqWrRmt_22 <= 6'h0;
      cntLkReqWrRmt_23 <= 6'h0;
      cntLkReqWrRmt_24 <= 6'h0;
      cntLkReqWrRmt_25 <= 6'h0;
      cntLkReqWrRmt_26 <= 6'h0;
      cntLkReqWrRmt_27 <= 6'h0;
      cntLkReqWrRmt_28 <= 6'h0;
      cntLkReqWrRmt_29 <= 6'h0;
      cntLkReqWrRmt_30 <= 6'h0;
      cntLkReqWrRmt_31 <= 6'h0;
      cntLkReqWrRmt_32 <= 6'h0;
      cntLkReqWrRmt_33 <= 6'h0;
      cntLkReqWrRmt_34 <= 6'h0;
      cntLkReqWrRmt_35 <= 6'h0;
      cntLkReqWrRmt_36 <= 6'h0;
      cntLkReqWrRmt_37 <= 6'h0;
      cntLkReqWrRmt_38 <= 6'h0;
      cntLkReqWrRmt_39 <= 6'h0;
      cntLkReqWrRmt_40 <= 6'h0;
      cntLkReqWrRmt_41 <= 6'h0;
      cntLkReqWrRmt_42 <= 6'h0;
      cntLkReqWrRmt_43 <= 6'h0;
      cntLkReqWrRmt_44 <= 6'h0;
      cntLkReqWrRmt_45 <= 6'h0;
      cntLkReqWrRmt_46 <= 6'h0;
      cntLkReqWrRmt_47 <= 6'h0;
      cntLkReqWrRmt_48 <= 6'h0;
      cntLkReqWrRmt_49 <= 6'h0;
      cntLkReqWrRmt_50 <= 6'h0;
      cntLkReqWrRmt_51 <= 6'h0;
      cntLkReqWrRmt_52 <= 6'h0;
      cntLkReqWrRmt_53 <= 6'h0;
      cntLkReqWrRmt_54 <= 6'h0;
      cntLkReqWrRmt_55 <= 6'h0;
      cntLkReqWrRmt_56 <= 6'h0;
      cntLkReqWrRmt_57 <= 6'h0;
      cntLkReqWrRmt_58 <= 6'h0;
      cntLkReqWrRmt_59 <= 6'h0;
      cntLkReqWrRmt_60 <= 6'h0;
      cntLkReqWrRmt_61 <= 6'h0;
      cntLkReqWrRmt_62 <= 6'h0;
      cntLkReqWrRmt_63 <= 6'h0;
      cntLkHoldWrLoc_0 <= 6'h0;
      cntLkHoldWrLoc_1 <= 6'h0;
      cntLkHoldWrLoc_2 <= 6'h0;
      cntLkHoldWrLoc_3 <= 6'h0;
      cntLkHoldWrLoc_4 <= 6'h0;
      cntLkHoldWrLoc_5 <= 6'h0;
      cntLkHoldWrLoc_6 <= 6'h0;
      cntLkHoldWrLoc_7 <= 6'h0;
      cntLkHoldWrLoc_8 <= 6'h0;
      cntLkHoldWrLoc_9 <= 6'h0;
      cntLkHoldWrLoc_10 <= 6'h0;
      cntLkHoldWrLoc_11 <= 6'h0;
      cntLkHoldWrLoc_12 <= 6'h0;
      cntLkHoldWrLoc_13 <= 6'h0;
      cntLkHoldWrLoc_14 <= 6'h0;
      cntLkHoldWrLoc_15 <= 6'h0;
      cntLkHoldWrLoc_16 <= 6'h0;
      cntLkHoldWrLoc_17 <= 6'h0;
      cntLkHoldWrLoc_18 <= 6'h0;
      cntLkHoldWrLoc_19 <= 6'h0;
      cntLkHoldWrLoc_20 <= 6'h0;
      cntLkHoldWrLoc_21 <= 6'h0;
      cntLkHoldWrLoc_22 <= 6'h0;
      cntLkHoldWrLoc_23 <= 6'h0;
      cntLkHoldWrLoc_24 <= 6'h0;
      cntLkHoldWrLoc_25 <= 6'h0;
      cntLkHoldWrLoc_26 <= 6'h0;
      cntLkHoldWrLoc_27 <= 6'h0;
      cntLkHoldWrLoc_28 <= 6'h0;
      cntLkHoldWrLoc_29 <= 6'h0;
      cntLkHoldWrLoc_30 <= 6'h0;
      cntLkHoldWrLoc_31 <= 6'h0;
      cntLkHoldWrLoc_32 <= 6'h0;
      cntLkHoldWrLoc_33 <= 6'h0;
      cntLkHoldWrLoc_34 <= 6'h0;
      cntLkHoldWrLoc_35 <= 6'h0;
      cntLkHoldWrLoc_36 <= 6'h0;
      cntLkHoldWrLoc_37 <= 6'h0;
      cntLkHoldWrLoc_38 <= 6'h0;
      cntLkHoldWrLoc_39 <= 6'h0;
      cntLkHoldWrLoc_40 <= 6'h0;
      cntLkHoldWrLoc_41 <= 6'h0;
      cntLkHoldWrLoc_42 <= 6'h0;
      cntLkHoldWrLoc_43 <= 6'h0;
      cntLkHoldWrLoc_44 <= 6'h0;
      cntLkHoldWrLoc_45 <= 6'h0;
      cntLkHoldWrLoc_46 <= 6'h0;
      cntLkHoldWrLoc_47 <= 6'h0;
      cntLkHoldWrLoc_48 <= 6'h0;
      cntLkHoldWrLoc_49 <= 6'h0;
      cntLkHoldWrLoc_50 <= 6'h0;
      cntLkHoldWrLoc_51 <= 6'h0;
      cntLkHoldWrLoc_52 <= 6'h0;
      cntLkHoldWrLoc_53 <= 6'h0;
      cntLkHoldWrLoc_54 <= 6'h0;
      cntLkHoldWrLoc_55 <= 6'h0;
      cntLkHoldWrLoc_56 <= 6'h0;
      cntLkHoldWrLoc_57 <= 6'h0;
      cntLkHoldWrLoc_58 <= 6'h0;
      cntLkHoldWrLoc_59 <= 6'h0;
      cntLkHoldWrLoc_60 <= 6'h0;
      cntLkHoldWrLoc_61 <= 6'h0;
      cntLkHoldWrLoc_62 <= 6'h0;
      cntLkHoldWrLoc_63 <= 6'h0;
      cntLkHoldWrRmt_0 <= 6'h0;
      cntLkHoldWrRmt_1 <= 6'h0;
      cntLkHoldWrRmt_2 <= 6'h0;
      cntLkHoldWrRmt_3 <= 6'h0;
      cntLkHoldWrRmt_4 <= 6'h0;
      cntLkHoldWrRmt_5 <= 6'h0;
      cntLkHoldWrRmt_6 <= 6'h0;
      cntLkHoldWrRmt_7 <= 6'h0;
      cntLkHoldWrRmt_8 <= 6'h0;
      cntLkHoldWrRmt_9 <= 6'h0;
      cntLkHoldWrRmt_10 <= 6'h0;
      cntLkHoldWrRmt_11 <= 6'h0;
      cntLkHoldWrRmt_12 <= 6'h0;
      cntLkHoldWrRmt_13 <= 6'h0;
      cntLkHoldWrRmt_14 <= 6'h0;
      cntLkHoldWrRmt_15 <= 6'h0;
      cntLkHoldWrRmt_16 <= 6'h0;
      cntLkHoldWrRmt_17 <= 6'h0;
      cntLkHoldWrRmt_18 <= 6'h0;
      cntLkHoldWrRmt_19 <= 6'h0;
      cntLkHoldWrRmt_20 <= 6'h0;
      cntLkHoldWrRmt_21 <= 6'h0;
      cntLkHoldWrRmt_22 <= 6'h0;
      cntLkHoldWrRmt_23 <= 6'h0;
      cntLkHoldWrRmt_24 <= 6'h0;
      cntLkHoldWrRmt_25 <= 6'h0;
      cntLkHoldWrRmt_26 <= 6'h0;
      cntLkHoldWrRmt_27 <= 6'h0;
      cntLkHoldWrRmt_28 <= 6'h0;
      cntLkHoldWrRmt_29 <= 6'h0;
      cntLkHoldWrRmt_30 <= 6'h0;
      cntLkHoldWrRmt_31 <= 6'h0;
      cntLkHoldWrRmt_32 <= 6'h0;
      cntLkHoldWrRmt_33 <= 6'h0;
      cntLkHoldWrRmt_34 <= 6'h0;
      cntLkHoldWrRmt_35 <= 6'h0;
      cntLkHoldWrRmt_36 <= 6'h0;
      cntLkHoldWrRmt_37 <= 6'h0;
      cntLkHoldWrRmt_38 <= 6'h0;
      cntLkHoldWrRmt_39 <= 6'h0;
      cntLkHoldWrRmt_40 <= 6'h0;
      cntLkHoldWrRmt_41 <= 6'h0;
      cntLkHoldWrRmt_42 <= 6'h0;
      cntLkHoldWrRmt_43 <= 6'h0;
      cntLkHoldWrRmt_44 <= 6'h0;
      cntLkHoldWrRmt_45 <= 6'h0;
      cntLkHoldWrRmt_46 <= 6'h0;
      cntLkHoldWrRmt_47 <= 6'h0;
      cntLkHoldWrRmt_48 <= 6'h0;
      cntLkHoldWrRmt_49 <= 6'h0;
      cntLkHoldWrRmt_50 <= 6'h0;
      cntLkHoldWrRmt_51 <= 6'h0;
      cntLkHoldWrRmt_52 <= 6'h0;
      cntLkHoldWrRmt_53 <= 6'h0;
      cntLkHoldWrRmt_54 <= 6'h0;
      cntLkHoldWrRmt_55 <= 6'h0;
      cntLkHoldWrRmt_56 <= 6'h0;
      cntLkHoldWrRmt_57 <= 6'h0;
      cntLkHoldWrRmt_58 <= 6'h0;
      cntLkHoldWrRmt_59 <= 6'h0;
      cntLkHoldWrRmt_60 <= 6'h0;
      cntLkHoldWrRmt_61 <= 6'h0;
      cntLkHoldWrRmt_62 <= 6'h0;
      cntLkHoldWrRmt_63 <= 6'h0;
      cntCmtReqLoc_0 <= 6'h0;
      cntCmtReqLoc_1 <= 6'h0;
      cntCmtReqLoc_2 <= 6'h0;
      cntCmtReqLoc_3 <= 6'h0;
      cntCmtReqLoc_4 <= 6'h0;
      cntCmtReqLoc_5 <= 6'h0;
      cntCmtReqLoc_6 <= 6'h0;
      cntCmtReqLoc_7 <= 6'h0;
      cntCmtReqLoc_8 <= 6'h0;
      cntCmtReqLoc_9 <= 6'h0;
      cntCmtReqLoc_10 <= 6'h0;
      cntCmtReqLoc_11 <= 6'h0;
      cntCmtReqLoc_12 <= 6'h0;
      cntCmtReqLoc_13 <= 6'h0;
      cntCmtReqLoc_14 <= 6'h0;
      cntCmtReqLoc_15 <= 6'h0;
      cntCmtReqLoc_16 <= 6'h0;
      cntCmtReqLoc_17 <= 6'h0;
      cntCmtReqLoc_18 <= 6'h0;
      cntCmtReqLoc_19 <= 6'h0;
      cntCmtReqLoc_20 <= 6'h0;
      cntCmtReqLoc_21 <= 6'h0;
      cntCmtReqLoc_22 <= 6'h0;
      cntCmtReqLoc_23 <= 6'h0;
      cntCmtReqLoc_24 <= 6'h0;
      cntCmtReqLoc_25 <= 6'h0;
      cntCmtReqLoc_26 <= 6'h0;
      cntCmtReqLoc_27 <= 6'h0;
      cntCmtReqLoc_28 <= 6'h0;
      cntCmtReqLoc_29 <= 6'h0;
      cntCmtReqLoc_30 <= 6'h0;
      cntCmtReqLoc_31 <= 6'h0;
      cntCmtReqLoc_32 <= 6'h0;
      cntCmtReqLoc_33 <= 6'h0;
      cntCmtReqLoc_34 <= 6'h0;
      cntCmtReqLoc_35 <= 6'h0;
      cntCmtReqLoc_36 <= 6'h0;
      cntCmtReqLoc_37 <= 6'h0;
      cntCmtReqLoc_38 <= 6'h0;
      cntCmtReqLoc_39 <= 6'h0;
      cntCmtReqLoc_40 <= 6'h0;
      cntCmtReqLoc_41 <= 6'h0;
      cntCmtReqLoc_42 <= 6'h0;
      cntCmtReqLoc_43 <= 6'h0;
      cntCmtReqLoc_44 <= 6'h0;
      cntCmtReqLoc_45 <= 6'h0;
      cntCmtReqLoc_46 <= 6'h0;
      cntCmtReqLoc_47 <= 6'h0;
      cntCmtReqLoc_48 <= 6'h0;
      cntCmtReqLoc_49 <= 6'h0;
      cntCmtReqLoc_50 <= 6'h0;
      cntCmtReqLoc_51 <= 6'h0;
      cntCmtReqLoc_52 <= 6'h0;
      cntCmtReqLoc_53 <= 6'h0;
      cntCmtReqLoc_54 <= 6'h0;
      cntCmtReqLoc_55 <= 6'h0;
      cntCmtReqLoc_56 <= 6'h0;
      cntCmtReqLoc_57 <= 6'h0;
      cntCmtReqLoc_58 <= 6'h0;
      cntCmtReqLoc_59 <= 6'h0;
      cntCmtReqLoc_60 <= 6'h0;
      cntCmtReqLoc_61 <= 6'h0;
      cntCmtReqLoc_62 <= 6'h0;
      cntCmtReqLoc_63 <= 6'h0;
      cntCmtReqRmt_0 <= 6'h0;
      cntCmtReqRmt_1 <= 6'h0;
      cntCmtReqRmt_2 <= 6'h0;
      cntCmtReqRmt_3 <= 6'h0;
      cntCmtReqRmt_4 <= 6'h0;
      cntCmtReqRmt_5 <= 6'h0;
      cntCmtReqRmt_6 <= 6'h0;
      cntCmtReqRmt_7 <= 6'h0;
      cntCmtReqRmt_8 <= 6'h0;
      cntCmtReqRmt_9 <= 6'h0;
      cntCmtReqRmt_10 <= 6'h0;
      cntCmtReqRmt_11 <= 6'h0;
      cntCmtReqRmt_12 <= 6'h0;
      cntCmtReqRmt_13 <= 6'h0;
      cntCmtReqRmt_14 <= 6'h0;
      cntCmtReqRmt_15 <= 6'h0;
      cntCmtReqRmt_16 <= 6'h0;
      cntCmtReqRmt_17 <= 6'h0;
      cntCmtReqRmt_18 <= 6'h0;
      cntCmtReqRmt_19 <= 6'h0;
      cntCmtReqRmt_20 <= 6'h0;
      cntCmtReqRmt_21 <= 6'h0;
      cntCmtReqRmt_22 <= 6'h0;
      cntCmtReqRmt_23 <= 6'h0;
      cntCmtReqRmt_24 <= 6'h0;
      cntCmtReqRmt_25 <= 6'h0;
      cntCmtReqRmt_26 <= 6'h0;
      cntCmtReqRmt_27 <= 6'h0;
      cntCmtReqRmt_28 <= 6'h0;
      cntCmtReqRmt_29 <= 6'h0;
      cntCmtReqRmt_30 <= 6'h0;
      cntCmtReqRmt_31 <= 6'h0;
      cntCmtReqRmt_32 <= 6'h0;
      cntCmtReqRmt_33 <= 6'h0;
      cntCmtReqRmt_34 <= 6'h0;
      cntCmtReqRmt_35 <= 6'h0;
      cntCmtReqRmt_36 <= 6'h0;
      cntCmtReqRmt_37 <= 6'h0;
      cntCmtReqRmt_38 <= 6'h0;
      cntCmtReqRmt_39 <= 6'h0;
      cntCmtReqRmt_40 <= 6'h0;
      cntCmtReqRmt_41 <= 6'h0;
      cntCmtReqRmt_42 <= 6'h0;
      cntCmtReqRmt_43 <= 6'h0;
      cntCmtReqRmt_44 <= 6'h0;
      cntCmtReqRmt_45 <= 6'h0;
      cntCmtReqRmt_46 <= 6'h0;
      cntCmtReqRmt_47 <= 6'h0;
      cntCmtReqRmt_48 <= 6'h0;
      cntCmtReqRmt_49 <= 6'h0;
      cntCmtReqRmt_50 <= 6'h0;
      cntCmtReqRmt_51 <= 6'h0;
      cntCmtReqRmt_52 <= 6'h0;
      cntCmtReqRmt_53 <= 6'h0;
      cntCmtReqRmt_54 <= 6'h0;
      cntCmtReqRmt_55 <= 6'h0;
      cntCmtReqRmt_56 <= 6'h0;
      cntCmtReqRmt_57 <= 6'h0;
      cntCmtReqRmt_58 <= 6'h0;
      cntCmtReqRmt_59 <= 6'h0;
      cntCmtReqRmt_60 <= 6'h0;
      cntCmtReqRmt_61 <= 6'h0;
      cntCmtReqRmt_62 <= 6'h0;
      cntCmtReqRmt_63 <= 6'h0;
      cntCmtRespLoc_0 <= 6'h0;
      cntCmtRespLoc_1 <= 6'h0;
      cntCmtRespLoc_2 <= 6'h0;
      cntCmtRespLoc_3 <= 6'h0;
      cntCmtRespLoc_4 <= 6'h0;
      cntCmtRespLoc_5 <= 6'h0;
      cntCmtRespLoc_6 <= 6'h0;
      cntCmtRespLoc_7 <= 6'h0;
      cntCmtRespLoc_8 <= 6'h0;
      cntCmtRespLoc_9 <= 6'h0;
      cntCmtRespLoc_10 <= 6'h0;
      cntCmtRespLoc_11 <= 6'h0;
      cntCmtRespLoc_12 <= 6'h0;
      cntCmtRespLoc_13 <= 6'h0;
      cntCmtRespLoc_14 <= 6'h0;
      cntCmtRespLoc_15 <= 6'h0;
      cntCmtRespLoc_16 <= 6'h0;
      cntCmtRespLoc_17 <= 6'h0;
      cntCmtRespLoc_18 <= 6'h0;
      cntCmtRespLoc_19 <= 6'h0;
      cntCmtRespLoc_20 <= 6'h0;
      cntCmtRespLoc_21 <= 6'h0;
      cntCmtRespLoc_22 <= 6'h0;
      cntCmtRespLoc_23 <= 6'h0;
      cntCmtRespLoc_24 <= 6'h0;
      cntCmtRespLoc_25 <= 6'h0;
      cntCmtRespLoc_26 <= 6'h0;
      cntCmtRespLoc_27 <= 6'h0;
      cntCmtRespLoc_28 <= 6'h0;
      cntCmtRespLoc_29 <= 6'h0;
      cntCmtRespLoc_30 <= 6'h0;
      cntCmtRespLoc_31 <= 6'h0;
      cntCmtRespLoc_32 <= 6'h0;
      cntCmtRespLoc_33 <= 6'h0;
      cntCmtRespLoc_34 <= 6'h0;
      cntCmtRespLoc_35 <= 6'h0;
      cntCmtRespLoc_36 <= 6'h0;
      cntCmtRespLoc_37 <= 6'h0;
      cntCmtRespLoc_38 <= 6'h0;
      cntCmtRespLoc_39 <= 6'h0;
      cntCmtRespLoc_40 <= 6'h0;
      cntCmtRespLoc_41 <= 6'h0;
      cntCmtRespLoc_42 <= 6'h0;
      cntCmtRespLoc_43 <= 6'h0;
      cntCmtRespLoc_44 <= 6'h0;
      cntCmtRespLoc_45 <= 6'h0;
      cntCmtRespLoc_46 <= 6'h0;
      cntCmtRespLoc_47 <= 6'h0;
      cntCmtRespLoc_48 <= 6'h0;
      cntCmtRespLoc_49 <= 6'h0;
      cntCmtRespLoc_50 <= 6'h0;
      cntCmtRespLoc_51 <= 6'h0;
      cntCmtRespLoc_52 <= 6'h0;
      cntCmtRespLoc_53 <= 6'h0;
      cntCmtRespLoc_54 <= 6'h0;
      cntCmtRespLoc_55 <= 6'h0;
      cntCmtRespLoc_56 <= 6'h0;
      cntCmtRespLoc_57 <= 6'h0;
      cntCmtRespLoc_58 <= 6'h0;
      cntCmtRespLoc_59 <= 6'h0;
      cntCmtRespLoc_60 <= 6'h0;
      cntCmtRespLoc_61 <= 6'h0;
      cntCmtRespLoc_62 <= 6'h0;
      cntCmtRespLoc_63 <= 6'h0;
      cntCmtRespRmt_0 <= 6'h0;
      cntCmtRespRmt_1 <= 6'h0;
      cntCmtRespRmt_2 <= 6'h0;
      cntCmtRespRmt_3 <= 6'h0;
      cntCmtRespRmt_4 <= 6'h0;
      cntCmtRespRmt_5 <= 6'h0;
      cntCmtRespRmt_6 <= 6'h0;
      cntCmtRespRmt_7 <= 6'h0;
      cntCmtRespRmt_8 <= 6'h0;
      cntCmtRespRmt_9 <= 6'h0;
      cntCmtRespRmt_10 <= 6'h0;
      cntCmtRespRmt_11 <= 6'h0;
      cntCmtRespRmt_12 <= 6'h0;
      cntCmtRespRmt_13 <= 6'h0;
      cntCmtRespRmt_14 <= 6'h0;
      cntCmtRespRmt_15 <= 6'h0;
      cntCmtRespRmt_16 <= 6'h0;
      cntCmtRespRmt_17 <= 6'h0;
      cntCmtRespRmt_18 <= 6'h0;
      cntCmtRespRmt_19 <= 6'h0;
      cntCmtRespRmt_20 <= 6'h0;
      cntCmtRespRmt_21 <= 6'h0;
      cntCmtRespRmt_22 <= 6'h0;
      cntCmtRespRmt_23 <= 6'h0;
      cntCmtRespRmt_24 <= 6'h0;
      cntCmtRespRmt_25 <= 6'h0;
      cntCmtRespRmt_26 <= 6'h0;
      cntCmtRespRmt_27 <= 6'h0;
      cntCmtRespRmt_28 <= 6'h0;
      cntCmtRespRmt_29 <= 6'h0;
      cntCmtRespRmt_30 <= 6'h0;
      cntCmtRespRmt_31 <= 6'h0;
      cntCmtRespRmt_32 <= 6'h0;
      cntCmtRespRmt_33 <= 6'h0;
      cntCmtRespRmt_34 <= 6'h0;
      cntCmtRespRmt_35 <= 6'h0;
      cntCmtRespRmt_36 <= 6'h0;
      cntCmtRespRmt_37 <= 6'h0;
      cntCmtRespRmt_38 <= 6'h0;
      cntCmtRespRmt_39 <= 6'h0;
      cntCmtRespRmt_40 <= 6'h0;
      cntCmtRespRmt_41 <= 6'h0;
      cntCmtRespRmt_42 <= 6'h0;
      cntCmtRespRmt_43 <= 6'h0;
      cntCmtRespRmt_44 <= 6'h0;
      cntCmtRespRmt_45 <= 6'h0;
      cntCmtRespRmt_46 <= 6'h0;
      cntCmtRespRmt_47 <= 6'h0;
      cntCmtRespRmt_48 <= 6'h0;
      cntCmtRespRmt_49 <= 6'h0;
      cntCmtRespRmt_50 <= 6'h0;
      cntCmtRespRmt_51 <= 6'h0;
      cntCmtRespRmt_52 <= 6'h0;
      cntCmtRespRmt_53 <= 6'h0;
      cntCmtRespRmt_54 <= 6'h0;
      cntCmtRespRmt_55 <= 6'h0;
      cntCmtRespRmt_56 <= 6'h0;
      cntCmtRespRmt_57 <= 6'h0;
      cntCmtRespRmt_58 <= 6'h0;
      cntCmtRespRmt_59 <= 6'h0;
      cntCmtRespRmt_60 <= 6'h0;
      cntCmtRespRmt_61 <= 6'h0;
      cntCmtRespRmt_62 <= 6'h0;
      cntCmtRespRmt_63 <= 6'h0;
      cntRlseReqLoc_0 <= 6'h0;
      cntRlseReqLoc_1 <= 6'h0;
      cntRlseReqLoc_2 <= 6'h0;
      cntRlseReqLoc_3 <= 6'h0;
      cntRlseReqLoc_4 <= 6'h0;
      cntRlseReqLoc_5 <= 6'h0;
      cntRlseReqLoc_6 <= 6'h0;
      cntRlseReqLoc_7 <= 6'h0;
      cntRlseReqLoc_8 <= 6'h0;
      cntRlseReqLoc_9 <= 6'h0;
      cntRlseReqLoc_10 <= 6'h0;
      cntRlseReqLoc_11 <= 6'h0;
      cntRlseReqLoc_12 <= 6'h0;
      cntRlseReqLoc_13 <= 6'h0;
      cntRlseReqLoc_14 <= 6'h0;
      cntRlseReqLoc_15 <= 6'h0;
      cntRlseReqLoc_16 <= 6'h0;
      cntRlseReqLoc_17 <= 6'h0;
      cntRlseReqLoc_18 <= 6'h0;
      cntRlseReqLoc_19 <= 6'h0;
      cntRlseReqLoc_20 <= 6'h0;
      cntRlseReqLoc_21 <= 6'h0;
      cntRlseReqLoc_22 <= 6'h0;
      cntRlseReqLoc_23 <= 6'h0;
      cntRlseReqLoc_24 <= 6'h0;
      cntRlseReqLoc_25 <= 6'h0;
      cntRlseReqLoc_26 <= 6'h0;
      cntRlseReqLoc_27 <= 6'h0;
      cntRlseReqLoc_28 <= 6'h0;
      cntRlseReqLoc_29 <= 6'h0;
      cntRlseReqLoc_30 <= 6'h0;
      cntRlseReqLoc_31 <= 6'h0;
      cntRlseReqLoc_32 <= 6'h0;
      cntRlseReqLoc_33 <= 6'h0;
      cntRlseReqLoc_34 <= 6'h0;
      cntRlseReqLoc_35 <= 6'h0;
      cntRlseReqLoc_36 <= 6'h0;
      cntRlseReqLoc_37 <= 6'h0;
      cntRlseReqLoc_38 <= 6'h0;
      cntRlseReqLoc_39 <= 6'h0;
      cntRlseReqLoc_40 <= 6'h0;
      cntRlseReqLoc_41 <= 6'h0;
      cntRlseReqLoc_42 <= 6'h0;
      cntRlseReqLoc_43 <= 6'h0;
      cntRlseReqLoc_44 <= 6'h0;
      cntRlseReqLoc_45 <= 6'h0;
      cntRlseReqLoc_46 <= 6'h0;
      cntRlseReqLoc_47 <= 6'h0;
      cntRlseReqLoc_48 <= 6'h0;
      cntRlseReqLoc_49 <= 6'h0;
      cntRlseReqLoc_50 <= 6'h0;
      cntRlseReqLoc_51 <= 6'h0;
      cntRlseReqLoc_52 <= 6'h0;
      cntRlseReqLoc_53 <= 6'h0;
      cntRlseReqLoc_54 <= 6'h0;
      cntRlseReqLoc_55 <= 6'h0;
      cntRlseReqLoc_56 <= 6'h0;
      cntRlseReqLoc_57 <= 6'h0;
      cntRlseReqLoc_58 <= 6'h0;
      cntRlseReqLoc_59 <= 6'h0;
      cntRlseReqLoc_60 <= 6'h0;
      cntRlseReqLoc_61 <= 6'h0;
      cntRlseReqLoc_62 <= 6'h0;
      cntRlseReqLoc_63 <= 6'h0;
      cntRlseReqRmt_0 <= 6'h0;
      cntRlseReqRmt_1 <= 6'h0;
      cntRlseReqRmt_2 <= 6'h0;
      cntRlseReqRmt_3 <= 6'h0;
      cntRlseReqRmt_4 <= 6'h0;
      cntRlseReqRmt_5 <= 6'h0;
      cntRlseReqRmt_6 <= 6'h0;
      cntRlseReqRmt_7 <= 6'h0;
      cntRlseReqRmt_8 <= 6'h0;
      cntRlseReqRmt_9 <= 6'h0;
      cntRlseReqRmt_10 <= 6'h0;
      cntRlseReqRmt_11 <= 6'h0;
      cntRlseReqRmt_12 <= 6'h0;
      cntRlseReqRmt_13 <= 6'h0;
      cntRlseReqRmt_14 <= 6'h0;
      cntRlseReqRmt_15 <= 6'h0;
      cntRlseReqRmt_16 <= 6'h0;
      cntRlseReqRmt_17 <= 6'h0;
      cntRlseReqRmt_18 <= 6'h0;
      cntRlseReqRmt_19 <= 6'h0;
      cntRlseReqRmt_20 <= 6'h0;
      cntRlseReqRmt_21 <= 6'h0;
      cntRlseReqRmt_22 <= 6'h0;
      cntRlseReqRmt_23 <= 6'h0;
      cntRlseReqRmt_24 <= 6'h0;
      cntRlseReqRmt_25 <= 6'h0;
      cntRlseReqRmt_26 <= 6'h0;
      cntRlseReqRmt_27 <= 6'h0;
      cntRlseReqRmt_28 <= 6'h0;
      cntRlseReqRmt_29 <= 6'h0;
      cntRlseReqRmt_30 <= 6'h0;
      cntRlseReqRmt_31 <= 6'h0;
      cntRlseReqRmt_32 <= 6'h0;
      cntRlseReqRmt_33 <= 6'h0;
      cntRlseReqRmt_34 <= 6'h0;
      cntRlseReqRmt_35 <= 6'h0;
      cntRlseReqRmt_36 <= 6'h0;
      cntRlseReqRmt_37 <= 6'h0;
      cntRlseReqRmt_38 <= 6'h0;
      cntRlseReqRmt_39 <= 6'h0;
      cntRlseReqRmt_40 <= 6'h0;
      cntRlseReqRmt_41 <= 6'h0;
      cntRlseReqRmt_42 <= 6'h0;
      cntRlseReqRmt_43 <= 6'h0;
      cntRlseReqRmt_44 <= 6'h0;
      cntRlseReqRmt_45 <= 6'h0;
      cntRlseReqRmt_46 <= 6'h0;
      cntRlseReqRmt_47 <= 6'h0;
      cntRlseReqRmt_48 <= 6'h0;
      cntRlseReqRmt_49 <= 6'h0;
      cntRlseReqRmt_50 <= 6'h0;
      cntRlseReqRmt_51 <= 6'h0;
      cntRlseReqRmt_52 <= 6'h0;
      cntRlseReqRmt_53 <= 6'h0;
      cntRlseReqRmt_54 <= 6'h0;
      cntRlseReqRmt_55 <= 6'h0;
      cntRlseReqRmt_56 <= 6'h0;
      cntRlseReqRmt_57 <= 6'h0;
      cntRlseReqRmt_58 <= 6'h0;
      cntRlseReqRmt_59 <= 6'h0;
      cntRlseReqRmt_60 <= 6'h0;
      cntRlseReqRmt_61 <= 6'h0;
      cntRlseReqRmt_62 <= 6'h0;
      cntRlseReqRmt_63 <= 6'h0;
      cntRlseReqWrLoc_0 <= 6'h0;
      cntRlseReqWrLoc_1 <= 6'h0;
      cntRlseReqWrLoc_2 <= 6'h0;
      cntRlseReqWrLoc_3 <= 6'h0;
      cntRlseReqWrLoc_4 <= 6'h0;
      cntRlseReqWrLoc_5 <= 6'h0;
      cntRlseReqWrLoc_6 <= 6'h0;
      cntRlseReqWrLoc_7 <= 6'h0;
      cntRlseReqWrLoc_8 <= 6'h0;
      cntRlseReqWrLoc_9 <= 6'h0;
      cntRlseReqWrLoc_10 <= 6'h0;
      cntRlseReqWrLoc_11 <= 6'h0;
      cntRlseReqWrLoc_12 <= 6'h0;
      cntRlseReqWrLoc_13 <= 6'h0;
      cntRlseReqWrLoc_14 <= 6'h0;
      cntRlseReqWrLoc_15 <= 6'h0;
      cntRlseReqWrLoc_16 <= 6'h0;
      cntRlseReqWrLoc_17 <= 6'h0;
      cntRlseReqWrLoc_18 <= 6'h0;
      cntRlseReqWrLoc_19 <= 6'h0;
      cntRlseReqWrLoc_20 <= 6'h0;
      cntRlseReqWrLoc_21 <= 6'h0;
      cntRlseReqWrLoc_22 <= 6'h0;
      cntRlseReqWrLoc_23 <= 6'h0;
      cntRlseReqWrLoc_24 <= 6'h0;
      cntRlseReqWrLoc_25 <= 6'h0;
      cntRlseReqWrLoc_26 <= 6'h0;
      cntRlseReqWrLoc_27 <= 6'h0;
      cntRlseReqWrLoc_28 <= 6'h0;
      cntRlseReqWrLoc_29 <= 6'h0;
      cntRlseReqWrLoc_30 <= 6'h0;
      cntRlseReqWrLoc_31 <= 6'h0;
      cntRlseReqWrLoc_32 <= 6'h0;
      cntRlseReqWrLoc_33 <= 6'h0;
      cntRlseReqWrLoc_34 <= 6'h0;
      cntRlseReqWrLoc_35 <= 6'h0;
      cntRlseReqWrLoc_36 <= 6'h0;
      cntRlseReqWrLoc_37 <= 6'h0;
      cntRlseReqWrLoc_38 <= 6'h0;
      cntRlseReqWrLoc_39 <= 6'h0;
      cntRlseReqWrLoc_40 <= 6'h0;
      cntRlseReqWrLoc_41 <= 6'h0;
      cntRlseReqWrLoc_42 <= 6'h0;
      cntRlseReqWrLoc_43 <= 6'h0;
      cntRlseReqWrLoc_44 <= 6'h0;
      cntRlseReqWrLoc_45 <= 6'h0;
      cntRlseReqWrLoc_46 <= 6'h0;
      cntRlseReqWrLoc_47 <= 6'h0;
      cntRlseReqWrLoc_48 <= 6'h0;
      cntRlseReqWrLoc_49 <= 6'h0;
      cntRlseReqWrLoc_50 <= 6'h0;
      cntRlseReqWrLoc_51 <= 6'h0;
      cntRlseReqWrLoc_52 <= 6'h0;
      cntRlseReqWrLoc_53 <= 6'h0;
      cntRlseReqWrLoc_54 <= 6'h0;
      cntRlseReqWrLoc_55 <= 6'h0;
      cntRlseReqWrLoc_56 <= 6'h0;
      cntRlseReqWrLoc_57 <= 6'h0;
      cntRlseReqWrLoc_58 <= 6'h0;
      cntRlseReqWrLoc_59 <= 6'h0;
      cntRlseReqWrLoc_60 <= 6'h0;
      cntRlseReqWrLoc_61 <= 6'h0;
      cntRlseReqWrLoc_62 <= 6'h0;
      cntRlseReqWrLoc_63 <= 6'h0;
      cntRlseReqWrRmt_0 <= 6'h0;
      cntRlseReqWrRmt_1 <= 6'h0;
      cntRlseReqWrRmt_2 <= 6'h0;
      cntRlseReqWrRmt_3 <= 6'h0;
      cntRlseReqWrRmt_4 <= 6'h0;
      cntRlseReqWrRmt_5 <= 6'h0;
      cntRlseReqWrRmt_6 <= 6'h0;
      cntRlseReqWrRmt_7 <= 6'h0;
      cntRlseReqWrRmt_8 <= 6'h0;
      cntRlseReqWrRmt_9 <= 6'h0;
      cntRlseReqWrRmt_10 <= 6'h0;
      cntRlseReqWrRmt_11 <= 6'h0;
      cntRlseReqWrRmt_12 <= 6'h0;
      cntRlseReqWrRmt_13 <= 6'h0;
      cntRlseReqWrRmt_14 <= 6'h0;
      cntRlseReqWrRmt_15 <= 6'h0;
      cntRlseReqWrRmt_16 <= 6'h0;
      cntRlseReqWrRmt_17 <= 6'h0;
      cntRlseReqWrRmt_18 <= 6'h0;
      cntRlseReqWrRmt_19 <= 6'h0;
      cntRlseReqWrRmt_20 <= 6'h0;
      cntRlseReqWrRmt_21 <= 6'h0;
      cntRlseReqWrRmt_22 <= 6'h0;
      cntRlseReqWrRmt_23 <= 6'h0;
      cntRlseReqWrRmt_24 <= 6'h0;
      cntRlseReqWrRmt_25 <= 6'h0;
      cntRlseReqWrRmt_26 <= 6'h0;
      cntRlseReqWrRmt_27 <= 6'h0;
      cntRlseReqWrRmt_28 <= 6'h0;
      cntRlseReqWrRmt_29 <= 6'h0;
      cntRlseReqWrRmt_30 <= 6'h0;
      cntRlseReqWrRmt_31 <= 6'h0;
      cntRlseReqWrRmt_32 <= 6'h0;
      cntRlseReqWrRmt_33 <= 6'h0;
      cntRlseReqWrRmt_34 <= 6'h0;
      cntRlseReqWrRmt_35 <= 6'h0;
      cntRlseReqWrRmt_36 <= 6'h0;
      cntRlseReqWrRmt_37 <= 6'h0;
      cntRlseReqWrRmt_38 <= 6'h0;
      cntRlseReqWrRmt_39 <= 6'h0;
      cntRlseReqWrRmt_40 <= 6'h0;
      cntRlseReqWrRmt_41 <= 6'h0;
      cntRlseReqWrRmt_42 <= 6'h0;
      cntRlseReqWrRmt_43 <= 6'h0;
      cntRlseReqWrRmt_44 <= 6'h0;
      cntRlseReqWrRmt_45 <= 6'h0;
      cntRlseReqWrRmt_46 <= 6'h0;
      cntRlseReqWrRmt_47 <= 6'h0;
      cntRlseReqWrRmt_48 <= 6'h0;
      cntRlseReqWrRmt_49 <= 6'h0;
      cntRlseReqWrRmt_50 <= 6'h0;
      cntRlseReqWrRmt_51 <= 6'h0;
      cntRlseReqWrRmt_52 <= 6'h0;
      cntRlseReqWrRmt_53 <= 6'h0;
      cntRlseReqWrRmt_54 <= 6'h0;
      cntRlseReqWrRmt_55 <= 6'h0;
      cntRlseReqWrRmt_56 <= 6'h0;
      cntRlseReqWrRmt_57 <= 6'h0;
      cntRlseReqWrRmt_58 <= 6'h0;
      cntRlseReqWrRmt_59 <= 6'h0;
      cntRlseReqWrRmt_60 <= 6'h0;
      cntRlseReqWrRmt_61 <= 6'h0;
      cntRlseReqWrRmt_62 <= 6'h0;
      cntRlseReqWrRmt_63 <= 6'h0;
      cntRlseRespLoc_0 <= 6'h0;
      cntRlseRespLoc_1 <= 6'h0;
      cntRlseRespLoc_2 <= 6'h0;
      cntRlseRespLoc_3 <= 6'h0;
      cntRlseRespLoc_4 <= 6'h0;
      cntRlseRespLoc_5 <= 6'h0;
      cntRlseRespLoc_6 <= 6'h0;
      cntRlseRespLoc_7 <= 6'h0;
      cntRlseRespLoc_8 <= 6'h0;
      cntRlseRespLoc_9 <= 6'h0;
      cntRlseRespLoc_10 <= 6'h0;
      cntRlseRespLoc_11 <= 6'h0;
      cntRlseRespLoc_12 <= 6'h0;
      cntRlseRespLoc_13 <= 6'h0;
      cntRlseRespLoc_14 <= 6'h0;
      cntRlseRespLoc_15 <= 6'h0;
      cntRlseRespLoc_16 <= 6'h0;
      cntRlseRespLoc_17 <= 6'h0;
      cntRlseRespLoc_18 <= 6'h0;
      cntRlseRespLoc_19 <= 6'h0;
      cntRlseRespLoc_20 <= 6'h0;
      cntRlseRespLoc_21 <= 6'h0;
      cntRlseRespLoc_22 <= 6'h0;
      cntRlseRespLoc_23 <= 6'h0;
      cntRlseRespLoc_24 <= 6'h0;
      cntRlseRespLoc_25 <= 6'h0;
      cntRlseRespLoc_26 <= 6'h0;
      cntRlseRespLoc_27 <= 6'h0;
      cntRlseRespLoc_28 <= 6'h0;
      cntRlseRespLoc_29 <= 6'h0;
      cntRlseRespLoc_30 <= 6'h0;
      cntRlseRespLoc_31 <= 6'h0;
      cntRlseRespLoc_32 <= 6'h0;
      cntRlseRespLoc_33 <= 6'h0;
      cntRlseRespLoc_34 <= 6'h0;
      cntRlseRespLoc_35 <= 6'h0;
      cntRlseRespLoc_36 <= 6'h0;
      cntRlseRespLoc_37 <= 6'h0;
      cntRlseRespLoc_38 <= 6'h0;
      cntRlseRespLoc_39 <= 6'h0;
      cntRlseRespLoc_40 <= 6'h0;
      cntRlseRespLoc_41 <= 6'h0;
      cntRlseRespLoc_42 <= 6'h0;
      cntRlseRespLoc_43 <= 6'h0;
      cntRlseRespLoc_44 <= 6'h0;
      cntRlseRespLoc_45 <= 6'h0;
      cntRlseRespLoc_46 <= 6'h0;
      cntRlseRespLoc_47 <= 6'h0;
      cntRlseRespLoc_48 <= 6'h0;
      cntRlseRespLoc_49 <= 6'h0;
      cntRlseRespLoc_50 <= 6'h0;
      cntRlseRespLoc_51 <= 6'h0;
      cntRlseRespLoc_52 <= 6'h0;
      cntRlseRespLoc_53 <= 6'h0;
      cntRlseRespLoc_54 <= 6'h0;
      cntRlseRespLoc_55 <= 6'h0;
      cntRlseRespLoc_56 <= 6'h0;
      cntRlseRespLoc_57 <= 6'h0;
      cntRlseRespLoc_58 <= 6'h0;
      cntRlseRespLoc_59 <= 6'h0;
      cntRlseRespLoc_60 <= 6'h0;
      cntRlseRespLoc_61 <= 6'h0;
      cntRlseRespLoc_62 <= 6'h0;
      cntRlseRespLoc_63 <= 6'h0;
      cntRlseRespRmt_0 <= 6'h0;
      cntRlseRespRmt_1 <= 6'h0;
      cntRlseRespRmt_2 <= 6'h0;
      cntRlseRespRmt_3 <= 6'h0;
      cntRlseRespRmt_4 <= 6'h0;
      cntRlseRespRmt_5 <= 6'h0;
      cntRlseRespRmt_6 <= 6'h0;
      cntRlseRespRmt_7 <= 6'h0;
      cntRlseRespRmt_8 <= 6'h0;
      cntRlseRespRmt_9 <= 6'h0;
      cntRlseRespRmt_10 <= 6'h0;
      cntRlseRespRmt_11 <= 6'h0;
      cntRlseRespRmt_12 <= 6'h0;
      cntRlseRespRmt_13 <= 6'h0;
      cntRlseRespRmt_14 <= 6'h0;
      cntRlseRespRmt_15 <= 6'h0;
      cntRlseRespRmt_16 <= 6'h0;
      cntRlseRespRmt_17 <= 6'h0;
      cntRlseRespRmt_18 <= 6'h0;
      cntRlseRespRmt_19 <= 6'h0;
      cntRlseRespRmt_20 <= 6'h0;
      cntRlseRespRmt_21 <= 6'h0;
      cntRlseRespRmt_22 <= 6'h0;
      cntRlseRespRmt_23 <= 6'h0;
      cntRlseRespRmt_24 <= 6'h0;
      cntRlseRespRmt_25 <= 6'h0;
      cntRlseRespRmt_26 <= 6'h0;
      cntRlseRespRmt_27 <= 6'h0;
      cntRlseRespRmt_28 <= 6'h0;
      cntRlseRespRmt_29 <= 6'h0;
      cntRlseRespRmt_30 <= 6'h0;
      cntRlseRespRmt_31 <= 6'h0;
      cntRlseRespRmt_32 <= 6'h0;
      cntRlseRespRmt_33 <= 6'h0;
      cntRlseRespRmt_34 <= 6'h0;
      cntRlseRespRmt_35 <= 6'h0;
      cntRlseRespRmt_36 <= 6'h0;
      cntRlseRespRmt_37 <= 6'h0;
      cntRlseRespRmt_38 <= 6'h0;
      cntRlseRespRmt_39 <= 6'h0;
      cntRlseRespRmt_40 <= 6'h0;
      cntRlseRespRmt_41 <= 6'h0;
      cntRlseRespRmt_42 <= 6'h0;
      cntRlseRespRmt_43 <= 6'h0;
      cntRlseRespRmt_44 <= 6'h0;
      cntRlseRespRmt_45 <= 6'h0;
      cntRlseRespRmt_46 <= 6'h0;
      cntRlseRespRmt_47 <= 6'h0;
      cntRlseRespRmt_48 <= 6'h0;
      cntRlseRespRmt_49 <= 6'h0;
      cntRlseRespRmt_50 <= 6'h0;
      cntRlseRespRmt_51 <= 6'h0;
      cntRlseRespRmt_52 <= 6'h0;
      cntRlseRespRmt_53 <= 6'h0;
      cntRlseRespRmt_54 <= 6'h0;
      cntRlseRespRmt_55 <= 6'h0;
      cntRlseRespRmt_56 <= 6'h0;
      cntRlseRespRmt_57 <= 6'h0;
      cntRlseRespRmt_58 <= 6'h0;
      cntRlseRespRmt_59 <= 6'h0;
      cntRlseRespRmt_60 <= 6'h0;
      cntRlseRespRmt_61 <= 6'h0;
      cntRlseRespRmt_62 <= 6'h0;
      cntRlseRespRmt_63 <= 6'h0;
      cntTimeOut_0 <= 24'h0;
      cntTimeOut_1 <= 24'h0;
      cntTimeOut_2 <= 24'h0;
      cntTimeOut_3 <= 24'h0;
      cntTimeOut_4 <= 24'h0;
      cntTimeOut_5 <= 24'h0;
      cntTimeOut_6 <= 24'h0;
      cntTimeOut_7 <= 24'h0;
      cntTimeOut_8 <= 24'h0;
      cntTimeOut_9 <= 24'h0;
      cntTimeOut_10 <= 24'h0;
      cntTimeOut_11 <= 24'h0;
      cntTimeOut_12 <= 24'h0;
      cntTimeOut_13 <= 24'h0;
      cntTimeOut_14 <= 24'h0;
      cntTimeOut_15 <= 24'h0;
      cntTimeOut_16 <= 24'h0;
      cntTimeOut_17 <= 24'h0;
      cntTimeOut_18 <= 24'h0;
      cntTimeOut_19 <= 24'h0;
      cntTimeOut_20 <= 24'h0;
      cntTimeOut_21 <= 24'h0;
      cntTimeOut_22 <= 24'h0;
      cntTimeOut_23 <= 24'h0;
      cntTimeOut_24 <= 24'h0;
      cntTimeOut_25 <= 24'h0;
      cntTimeOut_26 <= 24'h0;
      cntTimeOut_27 <= 24'h0;
      cntTimeOut_28 <= 24'h0;
      cntTimeOut_29 <= 24'h0;
      cntTimeOut_30 <= 24'h0;
      cntTimeOut_31 <= 24'h0;
      cntTimeOut_32 <= 24'h0;
      cntTimeOut_33 <= 24'h0;
      cntTimeOut_34 <= 24'h0;
      cntTimeOut_35 <= 24'h0;
      cntTimeOut_36 <= 24'h0;
      cntTimeOut_37 <= 24'h0;
      cntTimeOut_38 <= 24'h0;
      cntTimeOut_39 <= 24'h0;
      cntTimeOut_40 <= 24'h0;
      cntTimeOut_41 <= 24'h0;
      cntTimeOut_42 <= 24'h0;
      cntTimeOut_43 <= 24'h0;
      cntTimeOut_44 <= 24'h0;
      cntTimeOut_45 <= 24'h0;
      cntTimeOut_46 <= 24'h0;
      cntTimeOut_47 <= 24'h0;
      cntTimeOut_48 <= 24'h0;
      cntTimeOut_49 <= 24'h0;
      cntTimeOut_50 <= 24'h0;
      cntTimeOut_51 <= 24'h0;
      cntTimeOut_52 <= 24'h0;
      cntTimeOut_53 <= 24'h0;
      cntTimeOut_54 <= 24'h0;
      cntTimeOut_55 <= 24'h0;
      cntTimeOut_56 <= 24'h0;
      cntTimeOut_57 <= 24'h0;
      cntTimeOut_58 <= 24'h0;
      cntTimeOut_59 <= 24'h0;
      cntTimeOut_60 <= 24'h0;
      cntTimeOut_61 <= 24'h0;
      cntTimeOut_62 <= 24'h0;
      cntTimeOut_63 <= 24'h0;
      rTimeOut_0 <= 1'b0;
      rTimeOut_1 <= 1'b0;
      rTimeOut_2 <= 1'b0;
      rTimeOut_3 <= 1'b0;
      rTimeOut_4 <= 1'b0;
      rTimeOut_5 <= 1'b0;
      rTimeOut_6 <= 1'b0;
      rTimeOut_7 <= 1'b0;
      rTimeOut_8 <= 1'b0;
      rTimeOut_9 <= 1'b0;
      rTimeOut_10 <= 1'b0;
      rTimeOut_11 <= 1'b0;
      rTimeOut_12 <= 1'b0;
      rTimeOut_13 <= 1'b0;
      rTimeOut_14 <= 1'b0;
      rTimeOut_15 <= 1'b0;
      rTimeOut_16 <= 1'b0;
      rTimeOut_17 <= 1'b0;
      rTimeOut_18 <= 1'b0;
      rTimeOut_19 <= 1'b0;
      rTimeOut_20 <= 1'b0;
      rTimeOut_21 <= 1'b0;
      rTimeOut_22 <= 1'b0;
      rTimeOut_23 <= 1'b0;
      rTimeOut_24 <= 1'b0;
      rTimeOut_25 <= 1'b0;
      rTimeOut_26 <= 1'b0;
      rTimeOut_27 <= 1'b0;
      rTimeOut_28 <= 1'b0;
      rTimeOut_29 <= 1'b0;
      rTimeOut_30 <= 1'b0;
      rTimeOut_31 <= 1'b0;
      rTimeOut_32 <= 1'b0;
      rTimeOut_33 <= 1'b0;
      rTimeOut_34 <= 1'b0;
      rTimeOut_35 <= 1'b0;
      rTimeOut_36 <= 1'b0;
      rTimeOut_37 <= 1'b0;
      rTimeOut_38 <= 1'b0;
      rTimeOut_39 <= 1'b0;
      rTimeOut_40 <= 1'b0;
      rTimeOut_41 <= 1'b0;
      rTimeOut_42 <= 1'b0;
      rTimeOut_43 <= 1'b0;
      rTimeOut_44 <= 1'b0;
      rTimeOut_45 <= 1'b0;
      rTimeOut_46 <= 1'b0;
      rTimeOut_47 <= 1'b0;
      rTimeOut_48 <= 1'b0;
      rTimeOut_49 <= 1'b0;
      rTimeOut_50 <= 1'b0;
      rTimeOut_51 <= 1'b0;
      rTimeOut_52 <= 1'b0;
      rTimeOut_53 <= 1'b0;
      rTimeOut_54 <= 1'b0;
      rTimeOut_55 <= 1'b0;
      rTimeOut_56 <= 1'b0;
      rTimeOut_57 <= 1'b0;
      rTimeOut_58 <= 1'b0;
      rTimeOut_59 <= 1'b0;
      rTimeOut_60 <= 1'b0;
      rTimeOut_61 <= 1'b0;
      rTimeOut_62 <= 1'b0;
      rTimeOut_63 <= 1'b0;
      rAbort_0 <= 1'b0;
      rAbort_1 <= 1'b0;
      rAbort_2 <= 1'b0;
      rAbort_3 <= 1'b0;
      rAbort_4 <= 1'b0;
      rAbort_5 <= 1'b0;
      rAbort_6 <= 1'b0;
      rAbort_7 <= 1'b0;
      rAbort_8 <= 1'b0;
      rAbort_9 <= 1'b0;
      rAbort_10 <= 1'b0;
      rAbort_11 <= 1'b0;
      rAbort_12 <= 1'b0;
      rAbort_13 <= 1'b0;
      rAbort_14 <= 1'b0;
      rAbort_15 <= 1'b0;
      rAbort_16 <= 1'b0;
      rAbort_17 <= 1'b0;
      rAbort_18 <= 1'b0;
      rAbort_19 <= 1'b0;
      rAbort_20 <= 1'b0;
      rAbort_21 <= 1'b0;
      rAbort_22 <= 1'b0;
      rAbort_23 <= 1'b0;
      rAbort_24 <= 1'b0;
      rAbort_25 <= 1'b0;
      rAbort_26 <= 1'b0;
      rAbort_27 <= 1'b0;
      rAbort_28 <= 1'b0;
      rAbort_29 <= 1'b0;
      rAbort_30 <= 1'b0;
      rAbort_31 <= 1'b0;
      rAbort_32 <= 1'b0;
      rAbort_33 <= 1'b0;
      rAbort_34 <= 1'b0;
      rAbort_35 <= 1'b0;
      rAbort_36 <= 1'b0;
      rAbort_37 <= 1'b0;
      rAbort_38 <= 1'b0;
      rAbort_39 <= 1'b0;
      rAbort_40 <= 1'b0;
      rAbort_41 <= 1'b0;
      rAbort_42 <= 1'b0;
      rAbort_43 <= 1'b0;
      rAbort_44 <= 1'b0;
      rAbort_45 <= 1'b0;
      rAbort_46 <= 1'b0;
      rAbort_47 <= 1'b0;
      rAbort_48 <= 1'b0;
      rAbort_49 <= 1'b0;
      rAbort_50 <= 1'b0;
      rAbort_51 <= 1'b0;
      rAbort_52 <= 1'b0;
      rAbort_53 <= 1'b0;
      rAbort_54 <= 1'b0;
      rAbort_55 <= 1'b0;
      rAbort_56 <= 1'b0;
      rAbort_57 <= 1'b0;
      rAbort_58 <= 1'b0;
      rAbort_59 <= 1'b0;
      rAbort_60 <= 1'b0;
      rAbort_61 <= 1'b0;
      rAbort_62 <= 1'b0;
      rAbort_63 <= 1'b0;
      rReqDone_0 <= 1'b1;
      rReqDone_1 <= 1'b1;
      rReqDone_2 <= 1'b1;
      rReqDone_3 <= 1'b1;
      rReqDone_4 <= 1'b1;
      rReqDone_5 <= 1'b1;
      rReqDone_6 <= 1'b1;
      rReqDone_7 <= 1'b1;
      rReqDone_8 <= 1'b1;
      rReqDone_9 <= 1'b1;
      rReqDone_10 <= 1'b1;
      rReqDone_11 <= 1'b1;
      rReqDone_12 <= 1'b1;
      rReqDone_13 <= 1'b1;
      rReqDone_14 <= 1'b1;
      rReqDone_15 <= 1'b1;
      rReqDone_16 <= 1'b1;
      rReqDone_17 <= 1'b1;
      rReqDone_18 <= 1'b1;
      rReqDone_19 <= 1'b1;
      rReqDone_20 <= 1'b1;
      rReqDone_21 <= 1'b1;
      rReqDone_22 <= 1'b1;
      rReqDone_23 <= 1'b1;
      rReqDone_24 <= 1'b1;
      rReqDone_25 <= 1'b1;
      rReqDone_26 <= 1'b1;
      rReqDone_27 <= 1'b1;
      rReqDone_28 <= 1'b1;
      rReqDone_29 <= 1'b1;
      rReqDone_30 <= 1'b1;
      rReqDone_31 <= 1'b1;
      rReqDone_32 <= 1'b1;
      rReqDone_33 <= 1'b1;
      rReqDone_34 <= 1'b1;
      rReqDone_35 <= 1'b1;
      rReqDone_36 <= 1'b1;
      rReqDone_37 <= 1'b1;
      rReqDone_38 <= 1'b1;
      rReqDone_39 <= 1'b1;
      rReqDone_40 <= 1'b1;
      rReqDone_41 <= 1'b1;
      rReqDone_42 <= 1'b1;
      rReqDone_43 <= 1'b1;
      rReqDone_44 <= 1'b1;
      rReqDone_45 <= 1'b1;
      rReqDone_46 <= 1'b1;
      rReqDone_47 <= 1'b1;
      rReqDone_48 <= 1'b1;
      rReqDone_49 <= 1'b1;
      rReqDone_50 <= 1'b1;
      rReqDone_51 <= 1'b1;
      rReqDone_52 <= 1'b1;
      rReqDone_53 <= 1'b1;
      rReqDone_54 <= 1'b1;
      rReqDone_55 <= 1'b1;
      rReqDone_56 <= 1'b1;
      rReqDone_57 <= 1'b1;
      rReqDone_58 <= 1'b1;
      rReqDone_59 <= 1'b1;
      rReqDone_60 <= 1'b1;
      rReqDone_61 <= 1'b1;
      rReqDone_62 <= 1'b1;
      rReqDone_63 <= 1'b1;
      rRlseDone_0 <= 1'b1;
      rRlseDone_1 <= 1'b1;
      rRlseDone_2 <= 1'b1;
      rRlseDone_3 <= 1'b1;
      rRlseDone_4 <= 1'b1;
      rRlseDone_5 <= 1'b1;
      rRlseDone_6 <= 1'b1;
      rRlseDone_7 <= 1'b1;
      rRlseDone_8 <= 1'b1;
      rRlseDone_9 <= 1'b1;
      rRlseDone_10 <= 1'b1;
      rRlseDone_11 <= 1'b1;
      rRlseDone_12 <= 1'b1;
      rRlseDone_13 <= 1'b1;
      rRlseDone_14 <= 1'b1;
      rRlseDone_15 <= 1'b1;
      rRlseDone_16 <= 1'b1;
      rRlseDone_17 <= 1'b1;
      rRlseDone_18 <= 1'b1;
      rRlseDone_19 <= 1'b1;
      rRlseDone_20 <= 1'b1;
      rRlseDone_21 <= 1'b1;
      rRlseDone_22 <= 1'b1;
      rRlseDone_23 <= 1'b1;
      rRlseDone_24 <= 1'b1;
      rRlseDone_25 <= 1'b1;
      rRlseDone_26 <= 1'b1;
      rRlseDone_27 <= 1'b1;
      rRlseDone_28 <= 1'b1;
      rRlseDone_29 <= 1'b1;
      rRlseDone_30 <= 1'b1;
      rRlseDone_31 <= 1'b1;
      rRlseDone_32 <= 1'b1;
      rRlseDone_33 <= 1'b1;
      rRlseDone_34 <= 1'b1;
      rRlseDone_35 <= 1'b1;
      rRlseDone_36 <= 1'b1;
      rRlseDone_37 <= 1'b1;
      rRlseDone_38 <= 1'b1;
      rRlseDone_39 <= 1'b1;
      rRlseDone_40 <= 1'b1;
      rRlseDone_41 <= 1'b1;
      rRlseDone_42 <= 1'b1;
      rRlseDone_43 <= 1'b1;
      rRlseDone_44 <= 1'b1;
      rRlseDone_45 <= 1'b1;
      rRlseDone_46 <= 1'b1;
      rRlseDone_47 <= 1'b1;
      rRlseDone_48 <= 1'b1;
      rRlseDone_49 <= 1'b1;
      rRlseDone_50 <= 1'b1;
      rRlseDone_51 <= 1'b1;
      rRlseDone_52 <= 1'b1;
      rRlseDone_53 <= 1'b1;
      rRlseDone_54 <= 1'b1;
      rRlseDone_55 <= 1'b1;
      rRlseDone_56 <= 1'b1;
      rRlseDone_57 <= 1'b1;
      rRlseDone_58 <= 1'b1;
      rRlseDone_59 <= 1'b1;
      rRlseDone_60 <= 1'b1;
      rRlseDone_61 <= 1'b1;
      rRlseDone_62 <= 1'b1;
      rRlseDone_63 <= 1'b1;
      compLkReq_curTxnId <= 6'h0;
      _zz_compLkReq_txnMemRd_valid <= 1'b0;
      compLkReq_txnLen <= 6'h0;
      compLkReq_reqIdx <= 6'h0;
      compLkRespLoc_rFire <= 1'b0;
      compLkRespRmt_nBeat <= 8'h0;
      compLkRespRmt_rFire <= 1'b0;
      compTxnCmtLoc_curTxnId <= 6'h0;
      compTxnCmtLoc_nBeat <= 8'h0;
      compLkRlseLoc_curTxnId <= 6'h0;
      compLkRlseRmt_curTxnId <= 6'h0;
      compLkRlseRmt_nBeat <= 8'h0;
      compLoadTxn_curTxnId <= 6'h0;
      compLoadTxn_cntTxn <= 32'h0;
      compLoadTxn_rCmdAxiFire <= 1'b0;
      compLoadTxn_rTxnMemLd <= 1'b0;
      compLoadTxn_cntTxnWordInLine_value <= 3'b000;
      compLoadTxn_cntTxnWord_value <= 6'h0;
      compLkReq_stateReg <= compLkReq_enumDef_BOOT;
      compLkRespLoc_stateReg <= compLkRespLoc_enumDef_BOOT;
      compLkRespRmt_stateReg <= compLkRespRmt_enumDef_BOOT;
      compTxnCmtLoc_stateReg <= compTxnCmtLoc_enumDef_BOOT;
      compLkRlseLoc_stateReg <= compLkRlseLoc_enumDef_BOOT;
      compLkRlseRmt_stateReg <= compLkRlseRmt_enumDef_BOOT;
      compTimeOut_stateReg <= compTimeOut_enumDef_BOOT;
      compLoadTxn_stateReg <= compLoadTxn_enumDef_BOOT;
      clkCnt_stateReg <= clkCnt_enumDef_BOOT;
    end else begin
      if(streamArbiter_8_io_output_valid) begin
        streamArbiter_8_io_output_rValid <= 1'b1;
      end
      if(streamArbiter_8_io_output_s2mPipe_ready) begin
        streamArbiter_8_io_output_rValid <= 1'b0;
      end
      if(streamArbiter_8_io_output_s2mPipe_ready) begin
        streamArbiter_8_io_output_s2mPipe_rValid <= streamArbiter_8_io_output_s2mPipe_valid;
      end
      if(streamArbiter_9_io_output_valid) begin
        streamArbiter_9_io_output_rValid <= 1'b1;
      end
      if(streamArbiter_9_io_output_s2mPipe_ready) begin
        streamArbiter_9_io_output_rValid <= 1'b0;
      end
      if(streamArbiter_9_io_output_s2mPipe_ready) begin
        streamArbiter_9_io_output_s2mPipe_rValid <= streamArbiter_9_io_output_s2mPipe_valid;
      end
      if(compLkReq_txnMemRd_ready) begin
        _zz_compLkReq_txnMemRd_valid <= 1'b0;
      end
      if(compLkReq_txnMemRdCmd_ready) begin
        _zz_compLkReq_txnMemRd_valid <= compLkReq_txnMemRdCmd_valid;
      end
      compLkRespLoc_rFire <= io_lkRespLoc_fire_2;
      if(when_TxnManCS_l164) begin
        if(_zz_8[0]) begin
          rRlseDone_0 <= 1'b1;
        end
        if(_zz_8[1]) begin
          rRlseDone_1 <= 1'b1;
        end
        if(_zz_8[2]) begin
          rRlseDone_2 <= 1'b1;
        end
        if(_zz_8[3]) begin
          rRlseDone_3 <= 1'b1;
        end
        if(_zz_8[4]) begin
          rRlseDone_4 <= 1'b1;
        end
        if(_zz_8[5]) begin
          rRlseDone_5 <= 1'b1;
        end
        if(_zz_8[6]) begin
          rRlseDone_6 <= 1'b1;
        end
        if(_zz_8[7]) begin
          rRlseDone_7 <= 1'b1;
        end
        if(_zz_8[8]) begin
          rRlseDone_8 <= 1'b1;
        end
        if(_zz_8[9]) begin
          rRlseDone_9 <= 1'b1;
        end
        if(_zz_8[10]) begin
          rRlseDone_10 <= 1'b1;
        end
        if(_zz_8[11]) begin
          rRlseDone_11 <= 1'b1;
        end
        if(_zz_8[12]) begin
          rRlseDone_12 <= 1'b1;
        end
        if(_zz_8[13]) begin
          rRlseDone_13 <= 1'b1;
        end
        if(_zz_8[14]) begin
          rRlseDone_14 <= 1'b1;
        end
        if(_zz_8[15]) begin
          rRlseDone_15 <= 1'b1;
        end
        if(_zz_8[16]) begin
          rRlseDone_16 <= 1'b1;
        end
        if(_zz_8[17]) begin
          rRlseDone_17 <= 1'b1;
        end
        if(_zz_8[18]) begin
          rRlseDone_18 <= 1'b1;
        end
        if(_zz_8[19]) begin
          rRlseDone_19 <= 1'b1;
        end
        if(_zz_8[20]) begin
          rRlseDone_20 <= 1'b1;
        end
        if(_zz_8[21]) begin
          rRlseDone_21 <= 1'b1;
        end
        if(_zz_8[22]) begin
          rRlseDone_22 <= 1'b1;
        end
        if(_zz_8[23]) begin
          rRlseDone_23 <= 1'b1;
        end
        if(_zz_8[24]) begin
          rRlseDone_24 <= 1'b1;
        end
        if(_zz_8[25]) begin
          rRlseDone_25 <= 1'b1;
        end
        if(_zz_8[26]) begin
          rRlseDone_26 <= 1'b1;
        end
        if(_zz_8[27]) begin
          rRlseDone_27 <= 1'b1;
        end
        if(_zz_8[28]) begin
          rRlseDone_28 <= 1'b1;
        end
        if(_zz_8[29]) begin
          rRlseDone_29 <= 1'b1;
        end
        if(_zz_8[30]) begin
          rRlseDone_30 <= 1'b1;
        end
        if(_zz_8[31]) begin
          rRlseDone_31 <= 1'b1;
        end
        if(_zz_8[32]) begin
          rRlseDone_32 <= 1'b1;
        end
        if(_zz_8[33]) begin
          rRlseDone_33 <= 1'b1;
        end
        if(_zz_8[34]) begin
          rRlseDone_34 <= 1'b1;
        end
        if(_zz_8[35]) begin
          rRlseDone_35 <= 1'b1;
        end
        if(_zz_8[36]) begin
          rRlseDone_36 <= 1'b1;
        end
        if(_zz_8[37]) begin
          rRlseDone_37 <= 1'b1;
        end
        if(_zz_8[38]) begin
          rRlseDone_38 <= 1'b1;
        end
        if(_zz_8[39]) begin
          rRlseDone_39 <= 1'b1;
        end
        if(_zz_8[40]) begin
          rRlseDone_40 <= 1'b1;
        end
        if(_zz_8[41]) begin
          rRlseDone_41 <= 1'b1;
        end
        if(_zz_8[42]) begin
          rRlseDone_42 <= 1'b1;
        end
        if(_zz_8[43]) begin
          rRlseDone_43 <= 1'b1;
        end
        if(_zz_8[44]) begin
          rRlseDone_44 <= 1'b1;
        end
        if(_zz_8[45]) begin
          rRlseDone_45 <= 1'b1;
        end
        if(_zz_8[46]) begin
          rRlseDone_46 <= 1'b1;
        end
        if(_zz_8[47]) begin
          rRlseDone_47 <= 1'b1;
        end
        if(_zz_8[48]) begin
          rRlseDone_48 <= 1'b1;
        end
        if(_zz_8[49]) begin
          rRlseDone_49 <= 1'b1;
        end
        if(_zz_8[50]) begin
          rRlseDone_50 <= 1'b1;
        end
        if(_zz_8[51]) begin
          rRlseDone_51 <= 1'b1;
        end
        if(_zz_8[52]) begin
          rRlseDone_52 <= 1'b1;
        end
        if(_zz_8[53]) begin
          rRlseDone_53 <= 1'b1;
        end
        if(_zz_8[54]) begin
          rRlseDone_54 <= 1'b1;
        end
        if(_zz_8[55]) begin
          rRlseDone_55 <= 1'b1;
        end
        if(_zz_8[56]) begin
          rRlseDone_56 <= 1'b1;
        end
        if(_zz_8[57]) begin
          rRlseDone_57 <= 1'b1;
        end
        if(_zz_8[58]) begin
          rRlseDone_58 <= 1'b1;
        end
        if(_zz_8[59]) begin
          rRlseDone_59 <= 1'b1;
        end
        if(_zz_8[60]) begin
          rRlseDone_60 <= 1'b1;
        end
        if(_zz_8[61]) begin
          rRlseDone_61 <= 1'b1;
        end
        if(_zz_8[62]) begin
          rRlseDone_62 <= 1'b1;
        end
        if(_zz_8[63]) begin
          rRlseDone_63 <= 1'b1;
        end
        if(when_TxnManCS_l166) begin
          io_cntTxnAbt <= (io_cntTxnAbt + 32'h00000001);
        end else begin
          io_cntTxnCmt <= (io_cntTxnCmt + 32'h00000001);
        end
      end
      compLkRespRmt_rFire <= io_lkRespRmt_fire_2;
      if(when_TxnManCS_l259) begin
        if(_zz_12[0]) begin
          rRlseDone_0 <= 1'b1;
        end
        if(_zz_12[1]) begin
          rRlseDone_1 <= 1'b1;
        end
        if(_zz_12[2]) begin
          rRlseDone_2 <= 1'b1;
        end
        if(_zz_12[3]) begin
          rRlseDone_3 <= 1'b1;
        end
        if(_zz_12[4]) begin
          rRlseDone_4 <= 1'b1;
        end
        if(_zz_12[5]) begin
          rRlseDone_5 <= 1'b1;
        end
        if(_zz_12[6]) begin
          rRlseDone_6 <= 1'b1;
        end
        if(_zz_12[7]) begin
          rRlseDone_7 <= 1'b1;
        end
        if(_zz_12[8]) begin
          rRlseDone_8 <= 1'b1;
        end
        if(_zz_12[9]) begin
          rRlseDone_9 <= 1'b1;
        end
        if(_zz_12[10]) begin
          rRlseDone_10 <= 1'b1;
        end
        if(_zz_12[11]) begin
          rRlseDone_11 <= 1'b1;
        end
        if(_zz_12[12]) begin
          rRlseDone_12 <= 1'b1;
        end
        if(_zz_12[13]) begin
          rRlseDone_13 <= 1'b1;
        end
        if(_zz_12[14]) begin
          rRlseDone_14 <= 1'b1;
        end
        if(_zz_12[15]) begin
          rRlseDone_15 <= 1'b1;
        end
        if(_zz_12[16]) begin
          rRlseDone_16 <= 1'b1;
        end
        if(_zz_12[17]) begin
          rRlseDone_17 <= 1'b1;
        end
        if(_zz_12[18]) begin
          rRlseDone_18 <= 1'b1;
        end
        if(_zz_12[19]) begin
          rRlseDone_19 <= 1'b1;
        end
        if(_zz_12[20]) begin
          rRlseDone_20 <= 1'b1;
        end
        if(_zz_12[21]) begin
          rRlseDone_21 <= 1'b1;
        end
        if(_zz_12[22]) begin
          rRlseDone_22 <= 1'b1;
        end
        if(_zz_12[23]) begin
          rRlseDone_23 <= 1'b1;
        end
        if(_zz_12[24]) begin
          rRlseDone_24 <= 1'b1;
        end
        if(_zz_12[25]) begin
          rRlseDone_25 <= 1'b1;
        end
        if(_zz_12[26]) begin
          rRlseDone_26 <= 1'b1;
        end
        if(_zz_12[27]) begin
          rRlseDone_27 <= 1'b1;
        end
        if(_zz_12[28]) begin
          rRlseDone_28 <= 1'b1;
        end
        if(_zz_12[29]) begin
          rRlseDone_29 <= 1'b1;
        end
        if(_zz_12[30]) begin
          rRlseDone_30 <= 1'b1;
        end
        if(_zz_12[31]) begin
          rRlseDone_31 <= 1'b1;
        end
        if(_zz_12[32]) begin
          rRlseDone_32 <= 1'b1;
        end
        if(_zz_12[33]) begin
          rRlseDone_33 <= 1'b1;
        end
        if(_zz_12[34]) begin
          rRlseDone_34 <= 1'b1;
        end
        if(_zz_12[35]) begin
          rRlseDone_35 <= 1'b1;
        end
        if(_zz_12[36]) begin
          rRlseDone_36 <= 1'b1;
        end
        if(_zz_12[37]) begin
          rRlseDone_37 <= 1'b1;
        end
        if(_zz_12[38]) begin
          rRlseDone_38 <= 1'b1;
        end
        if(_zz_12[39]) begin
          rRlseDone_39 <= 1'b1;
        end
        if(_zz_12[40]) begin
          rRlseDone_40 <= 1'b1;
        end
        if(_zz_12[41]) begin
          rRlseDone_41 <= 1'b1;
        end
        if(_zz_12[42]) begin
          rRlseDone_42 <= 1'b1;
        end
        if(_zz_12[43]) begin
          rRlseDone_43 <= 1'b1;
        end
        if(_zz_12[44]) begin
          rRlseDone_44 <= 1'b1;
        end
        if(_zz_12[45]) begin
          rRlseDone_45 <= 1'b1;
        end
        if(_zz_12[46]) begin
          rRlseDone_46 <= 1'b1;
        end
        if(_zz_12[47]) begin
          rRlseDone_47 <= 1'b1;
        end
        if(_zz_12[48]) begin
          rRlseDone_48 <= 1'b1;
        end
        if(_zz_12[49]) begin
          rRlseDone_49 <= 1'b1;
        end
        if(_zz_12[50]) begin
          rRlseDone_50 <= 1'b1;
        end
        if(_zz_12[51]) begin
          rRlseDone_51 <= 1'b1;
        end
        if(_zz_12[52]) begin
          rRlseDone_52 <= 1'b1;
        end
        if(_zz_12[53]) begin
          rRlseDone_53 <= 1'b1;
        end
        if(_zz_12[54]) begin
          rRlseDone_54 <= 1'b1;
        end
        if(_zz_12[55]) begin
          rRlseDone_55 <= 1'b1;
        end
        if(_zz_12[56]) begin
          rRlseDone_56 <= 1'b1;
        end
        if(_zz_12[57]) begin
          rRlseDone_57 <= 1'b1;
        end
        if(_zz_12[58]) begin
          rRlseDone_58 <= 1'b1;
        end
        if(_zz_12[59]) begin
          rRlseDone_59 <= 1'b1;
        end
        if(_zz_12[60]) begin
          rRlseDone_60 <= 1'b1;
        end
        if(_zz_12[61]) begin
          rRlseDone_61 <= 1'b1;
        end
        if(_zz_12[62]) begin
          rRlseDone_62 <= 1'b1;
        end
        if(_zz_12[63]) begin
          rRlseDone_63 <= 1'b1;
        end
        if(when_TxnManCS_l261) begin
          io_cntTxnAbt <= (io_cntTxnAbt + 32'h00000001);
        end else begin
          io_cntTxnCmt <= (io_cntTxnCmt + 32'h00000001);
        end
      end
      if(compAxiResp_rAxiBFire) begin
        if(_zz_13[0]) begin
          cntCmtRespLoc_0 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[1]) begin
          cntCmtRespLoc_1 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[2]) begin
          cntCmtRespLoc_2 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[3]) begin
          cntCmtRespLoc_3 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[4]) begin
          cntCmtRespLoc_4 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[5]) begin
          cntCmtRespLoc_5 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[6]) begin
          cntCmtRespLoc_6 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[7]) begin
          cntCmtRespLoc_7 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[8]) begin
          cntCmtRespLoc_8 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[9]) begin
          cntCmtRespLoc_9 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[10]) begin
          cntCmtRespLoc_10 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[11]) begin
          cntCmtRespLoc_11 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[12]) begin
          cntCmtRespLoc_12 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[13]) begin
          cntCmtRespLoc_13 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[14]) begin
          cntCmtRespLoc_14 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[15]) begin
          cntCmtRespLoc_15 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[16]) begin
          cntCmtRespLoc_16 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[17]) begin
          cntCmtRespLoc_17 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[18]) begin
          cntCmtRespLoc_18 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[19]) begin
          cntCmtRespLoc_19 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[20]) begin
          cntCmtRespLoc_20 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[21]) begin
          cntCmtRespLoc_21 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[22]) begin
          cntCmtRespLoc_22 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[23]) begin
          cntCmtRespLoc_23 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[24]) begin
          cntCmtRespLoc_24 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[25]) begin
          cntCmtRespLoc_25 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[26]) begin
          cntCmtRespLoc_26 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[27]) begin
          cntCmtRespLoc_27 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[28]) begin
          cntCmtRespLoc_28 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[29]) begin
          cntCmtRespLoc_29 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[30]) begin
          cntCmtRespLoc_30 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[31]) begin
          cntCmtRespLoc_31 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[32]) begin
          cntCmtRespLoc_32 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[33]) begin
          cntCmtRespLoc_33 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[34]) begin
          cntCmtRespLoc_34 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[35]) begin
          cntCmtRespLoc_35 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[36]) begin
          cntCmtRespLoc_36 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[37]) begin
          cntCmtRespLoc_37 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[38]) begin
          cntCmtRespLoc_38 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[39]) begin
          cntCmtRespLoc_39 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[40]) begin
          cntCmtRespLoc_40 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[41]) begin
          cntCmtRespLoc_41 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[42]) begin
          cntCmtRespLoc_42 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[43]) begin
          cntCmtRespLoc_43 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[44]) begin
          cntCmtRespLoc_44 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[45]) begin
          cntCmtRespLoc_45 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[46]) begin
          cntCmtRespLoc_46 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[47]) begin
          cntCmtRespLoc_47 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[48]) begin
          cntCmtRespLoc_48 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[49]) begin
          cntCmtRespLoc_49 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[50]) begin
          cntCmtRespLoc_50 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[51]) begin
          cntCmtRespLoc_51 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[52]) begin
          cntCmtRespLoc_52 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[53]) begin
          cntCmtRespLoc_53 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[54]) begin
          cntCmtRespLoc_54 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[55]) begin
          cntCmtRespLoc_55 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[56]) begin
          cntCmtRespLoc_56 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[57]) begin
          cntCmtRespLoc_57 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[58]) begin
          cntCmtRespLoc_58 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[59]) begin
          cntCmtRespLoc_59 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[60]) begin
          cntCmtRespLoc_60 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[61]) begin
          cntCmtRespLoc_61 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[62]) begin
          cntCmtRespLoc_62 <= _zz_cntCmtRespLoc_0;
        end
        if(_zz_13[63]) begin
          cntCmtRespLoc_63 <= _zz_cntCmtRespLoc_0;
        end
      end
      compLoadTxn_rCmdAxiFire <= io_cmdAxi_r_fire_1;
      compLoadTxn_cntTxnWordInLine_value <= compLoadTxn_cntTxnWordInLine_valueNext;
      compLoadTxn_cntTxnWord_value <= compLoadTxn_cntTxnWord_valueNext;
      if(when_TxnManCS_l672) begin
        io_done <= 1'b1;
      end
      compLkReq_stateReg <= compLkReq_stateNext;
      case(compLkReq_stateReg)
        compLkReq_enumDef_CS_TXN : begin
          if(_zz_81) begin
            compLkReq_curTxnId <= compLkReq_rIdxTxn2Start;
          end
          if(compLkReq_txnMemRd_fire) begin
            compLkReq_txnLen <= _zz_compLkReq_txnLen[5 : 0];
          end
        end
        compLkReq_enumDef_RD_TXN : begin
          if(compLkReq_lkReqFire) begin
            compLkReq_reqIdx <= (compLkReq_reqIdx + 6'h01);
            case(compLkReq_isLocal)
              1'b1 : begin
                if(_zz_82[0]) begin
                  cntLkReqLoc_0 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[1]) begin
                  cntLkReqLoc_1 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[2]) begin
                  cntLkReqLoc_2 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[3]) begin
                  cntLkReqLoc_3 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[4]) begin
                  cntLkReqLoc_4 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[5]) begin
                  cntLkReqLoc_5 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[6]) begin
                  cntLkReqLoc_6 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[7]) begin
                  cntLkReqLoc_7 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[8]) begin
                  cntLkReqLoc_8 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[9]) begin
                  cntLkReqLoc_9 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[10]) begin
                  cntLkReqLoc_10 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[11]) begin
                  cntLkReqLoc_11 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[12]) begin
                  cntLkReqLoc_12 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[13]) begin
                  cntLkReqLoc_13 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[14]) begin
                  cntLkReqLoc_14 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[15]) begin
                  cntLkReqLoc_15 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[16]) begin
                  cntLkReqLoc_16 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[17]) begin
                  cntLkReqLoc_17 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[18]) begin
                  cntLkReqLoc_18 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[19]) begin
                  cntLkReqLoc_19 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[20]) begin
                  cntLkReqLoc_20 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[21]) begin
                  cntLkReqLoc_21 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[22]) begin
                  cntLkReqLoc_22 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[23]) begin
                  cntLkReqLoc_23 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[24]) begin
                  cntLkReqLoc_24 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[25]) begin
                  cntLkReqLoc_25 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[26]) begin
                  cntLkReqLoc_26 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[27]) begin
                  cntLkReqLoc_27 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[28]) begin
                  cntLkReqLoc_28 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[29]) begin
                  cntLkReqLoc_29 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[30]) begin
                  cntLkReqLoc_30 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[31]) begin
                  cntLkReqLoc_31 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[32]) begin
                  cntLkReqLoc_32 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[33]) begin
                  cntLkReqLoc_33 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[34]) begin
                  cntLkReqLoc_34 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[35]) begin
                  cntLkReqLoc_35 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[36]) begin
                  cntLkReqLoc_36 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[37]) begin
                  cntLkReqLoc_37 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[38]) begin
                  cntLkReqLoc_38 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[39]) begin
                  cntLkReqLoc_39 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[40]) begin
                  cntLkReqLoc_40 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[41]) begin
                  cntLkReqLoc_41 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[42]) begin
                  cntLkReqLoc_42 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[43]) begin
                  cntLkReqLoc_43 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[44]) begin
                  cntLkReqLoc_44 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[45]) begin
                  cntLkReqLoc_45 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[46]) begin
                  cntLkReqLoc_46 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[47]) begin
                  cntLkReqLoc_47 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[48]) begin
                  cntLkReqLoc_48 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[49]) begin
                  cntLkReqLoc_49 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[50]) begin
                  cntLkReqLoc_50 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[51]) begin
                  cntLkReqLoc_51 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[52]) begin
                  cntLkReqLoc_52 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[53]) begin
                  cntLkReqLoc_53 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[54]) begin
                  cntLkReqLoc_54 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[55]) begin
                  cntLkReqLoc_55 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[56]) begin
                  cntLkReqLoc_56 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[57]) begin
                  cntLkReqLoc_57 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[58]) begin
                  cntLkReqLoc_58 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[59]) begin
                  cntLkReqLoc_59 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[60]) begin
                  cntLkReqLoc_60 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[61]) begin
                  cntLkReqLoc_61 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[62]) begin
                  cntLkReqLoc_62 <= _zz_cntLkReqLoc_0;
                end
                if(_zz_82[63]) begin
                  cntLkReqLoc_63 <= _zz_cntLkReqLoc_0;
                end
                io_cntLockLoc <= (io_cntLockLoc + 32'h00000001);
              end
              default : begin
                if(_zz_83[0]) begin
                  cntLkReqRmt_0 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[1]) begin
                  cntLkReqRmt_1 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[2]) begin
                  cntLkReqRmt_2 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[3]) begin
                  cntLkReqRmt_3 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[4]) begin
                  cntLkReqRmt_4 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[5]) begin
                  cntLkReqRmt_5 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[6]) begin
                  cntLkReqRmt_6 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[7]) begin
                  cntLkReqRmt_7 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[8]) begin
                  cntLkReqRmt_8 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[9]) begin
                  cntLkReqRmt_9 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[10]) begin
                  cntLkReqRmt_10 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[11]) begin
                  cntLkReqRmt_11 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[12]) begin
                  cntLkReqRmt_12 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[13]) begin
                  cntLkReqRmt_13 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[14]) begin
                  cntLkReqRmt_14 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[15]) begin
                  cntLkReqRmt_15 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[16]) begin
                  cntLkReqRmt_16 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[17]) begin
                  cntLkReqRmt_17 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[18]) begin
                  cntLkReqRmt_18 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[19]) begin
                  cntLkReqRmt_19 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[20]) begin
                  cntLkReqRmt_20 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[21]) begin
                  cntLkReqRmt_21 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[22]) begin
                  cntLkReqRmt_22 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[23]) begin
                  cntLkReqRmt_23 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[24]) begin
                  cntLkReqRmt_24 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[25]) begin
                  cntLkReqRmt_25 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[26]) begin
                  cntLkReqRmt_26 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[27]) begin
                  cntLkReqRmt_27 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[28]) begin
                  cntLkReqRmt_28 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[29]) begin
                  cntLkReqRmt_29 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[30]) begin
                  cntLkReqRmt_30 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[31]) begin
                  cntLkReqRmt_31 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[32]) begin
                  cntLkReqRmt_32 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[33]) begin
                  cntLkReqRmt_33 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[34]) begin
                  cntLkReqRmt_34 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[35]) begin
                  cntLkReqRmt_35 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[36]) begin
                  cntLkReqRmt_36 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[37]) begin
                  cntLkReqRmt_37 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[38]) begin
                  cntLkReqRmt_38 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[39]) begin
                  cntLkReqRmt_39 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[40]) begin
                  cntLkReqRmt_40 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[41]) begin
                  cntLkReqRmt_41 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[42]) begin
                  cntLkReqRmt_42 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[43]) begin
                  cntLkReqRmt_43 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[44]) begin
                  cntLkReqRmt_44 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[45]) begin
                  cntLkReqRmt_45 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[46]) begin
                  cntLkReqRmt_46 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[47]) begin
                  cntLkReqRmt_47 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[48]) begin
                  cntLkReqRmt_48 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[49]) begin
                  cntLkReqRmt_49 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[50]) begin
                  cntLkReqRmt_50 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[51]) begin
                  cntLkReqRmt_51 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[52]) begin
                  cntLkReqRmt_52 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[53]) begin
                  cntLkReqRmt_53 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[54]) begin
                  cntLkReqRmt_54 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[55]) begin
                  cntLkReqRmt_55 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[56]) begin
                  cntLkReqRmt_56 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[57]) begin
                  cntLkReqRmt_57 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[58]) begin
                  cntLkReqRmt_58 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[59]) begin
                  cntLkReqRmt_59 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[60]) begin
                  cntLkReqRmt_60 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[61]) begin
                  cntLkReqRmt_61 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[62]) begin
                  cntLkReqRmt_62 <= _zz_cntLkReqRmt_0;
                end
                if(_zz_83[63]) begin
                  cntLkReqRmt_63 <= _zz_cntLkReqRmt_0;
                end
                io_cntLockRmt <= (io_cntLockRmt + 32'h00000001);
              end
            endcase
            if(when_TxnManCS_l106) begin
              case(compLkReq_isLocal)
                1'b1 : begin
                  if(_zz_84[0]) begin
                    cntLkReqWrLoc_0 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[1]) begin
                    cntLkReqWrLoc_1 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[2]) begin
                    cntLkReqWrLoc_2 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[3]) begin
                    cntLkReqWrLoc_3 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[4]) begin
                    cntLkReqWrLoc_4 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[5]) begin
                    cntLkReqWrLoc_5 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[6]) begin
                    cntLkReqWrLoc_6 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[7]) begin
                    cntLkReqWrLoc_7 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[8]) begin
                    cntLkReqWrLoc_8 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[9]) begin
                    cntLkReqWrLoc_9 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[10]) begin
                    cntLkReqWrLoc_10 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[11]) begin
                    cntLkReqWrLoc_11 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[12]) begin
                    cntLkReqWrLoc_12 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[13]) begin
                    cntLkReqWrLoc_13 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[14]) begin
                    cntLkReqWrLoc_14 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[15]) begin
                    cntLkReqWrLoc_15 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[16]) begin
                    cntLkReqWrLoc_16 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[17]) begin
                    cntLkReqWrLoc_17 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[18]) begin
                    cntLkReqWrLoc_18 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[19]) begin
                    cntLkReqWrLoc_19 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[20]) begin
                    cntLkReqWrLoc_20 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[21]) begin
                    cntLkReqWrLoc_21 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[22]) begin
                    cntLkReqWrLoc_22 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[23]) begin
                    cntLkReqWrLoc_23 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[24]) begin
                    cntLkReqWrLoc_24 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[25]) begin
                    cntLkReqWrLoc_25 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[26]) begin
                    cntLkReqWrLoc_26 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[27]) begin
                    cntLkReqWrLoc_27 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[28]) begin
                    cntLkReqWrLoc_28 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[29]) begin
                    cntLkReqWrLoc_29 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[30]) begin
                    cntLkReqWrLoc_30 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[31]) begin
                    cntLkReqWrLoc_31 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[32]) begin
                    cntLkReqWrLoc_32 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[33]) begin
                    cntLkReqWrLoc_33 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[34]) begin
                    cntLkReqWrLoc_34 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[35]) begin
                    cntLkReqWrLoc_35 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[36]) begin
                    cntLkReqWrLoc_36 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[37]) begin
                    cntLkReqWrLoc_37 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[38]) begin
                    cntLkReqWrLoc_38 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[39]) begin
                    cntLkReqWrLoc_39 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[40]) begin
                    cntLkReqWrLoc_40 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[41]) begin
                    cntLkReqWrLoc_41 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[42]) begin
                    cntLkReqWrLoc_42 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[43]) begin
                    cntLkReqWrLoc_43 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[44]) begin
                    cntLkReqWrLoc_44 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[45]) begin
                    cntLkReqWrLoc_45 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[46]) begin
                    cntLkReqWrLoc_46 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[47]) begin
                    cntLkReqWrLoc_47 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[48]) begin
                    cntLkReqWrLoc_48 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[49]) begin
                    cntLkReqWrLoc_49 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[50]) begin
                    cntLkReqWrLoc_50 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[51]) begin
                    cntLkReqWrLoc_51 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[52]) begin
                    cntLkReqWrLoc_52 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[53]) begin
                    cntLkReqWrLoc_53 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[54]) begin
                    cntLkReqWrLoc_54 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[55]) begin
                    cntLkReqWrLoc_55 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[56]) begin
                    cntLkReqWrLoc_56 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[57]) begin
                    cntLkReqWrLoc_57 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[58]) begin
                    cntLkReqWrLoc_58 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[59]) begin
                    cntLkReqWrLoc_59 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[60]) begin
                    cntLkReqWrLoc_60 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[61]) begin
                    cntLkReqWrLoc_61 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[62]) begin
                    cntLkReqWrLoc_62 <= _zz_cntLkReqWrLoc_0_1;
                  end
                  if(_zz_84[63]) begin
                    cntLkReqWrLoc_63 <= _zz_cntLkReqWrLoc_0_1;
                  end
                end
                default : begin
                  if(_zz_85[0]) begin
                    cntLkReqWrRmt_0 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[1]) begin
                    cntLkReqWrRmt_1 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[2]) begin
                    cntLkReqWrRmt_2 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[3]) begin
                    cntLkReqWrRmt_3 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[4]) begin
                    cntLkReqWrRmt_4 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[5]) begin
                    cntLkReqWrRmt_5 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[6]) begin
                    cntLkReqWrRmt_6 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[7]) begin
                    cntLkReqWrRmt_7 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[8]) begin
                    cntLkReqWrRmt_8 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[9]) begin
                    cntLkReqWrRmt_9 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[10]) begin
                    cntLkReqWrRmt_10 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[11]) begin
                    cntLkReqWrRmt_11 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[12]) begin
                    cntLkReqWrRmt_12 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[13]) begin
                    cntLkReqWrRmt_13 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[14]) begin
                    cntLkReqWrRmt_14 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[15]) begin
                    cntLkReqWrRmt_15 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[16]) begin
                    cntLkReqWrRmt_16 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[17]) begin
                    cntLkReqWrRmt_17 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[18]) begin
                    cntLkReqWrRmt_18 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[19]) begin
                    cntLkReqWrRmt_19 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[20]) begin
                    cntLkReqWrRmt_20 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[21]) begin
                    cntLkReqWrRmt_21 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[22]) begin
                    cntLkReqWrRmt_22 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[23]) begin
                    cntLkReqWrRmt_23 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[24]) begin
                    cntLkReqWrRmt_24 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[25]) begin
                    cntLkReqWrRmt_25 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[26]) begin
                    cntLkReqWrRmt_26 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[27]) begin
                    cntLkReqWrRmt_27 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[28]) begin
                    cntLkReqWrRmt_28 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[29]) begin
                    cntLkReqWrRmt_29 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[30]) begin
                    cntLkReqWrRmt_30 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[31]) begin
                    cntLkReqWrRmt_31 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[32]) begin
                    cntLkReqWrRmt_32 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[33]) begin
                    cntLkReqWrRmt_33 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[34]) begin
                    cntLkReqWrRmt_34 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[35]) begin
                    cntLkReqWrRmt_35 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[36]) begin
                    cntLkReqWrRmt_36 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[37]) begin
                    cntLkReqWrRmt_37 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[38]) begin
                    cntLkReqWrRmt_38 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[39]) begin
                    cntLkReqWrRmt_39 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[40]) begin
                    cntLkReqWrRmt_40 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[41]) begin
                    cntLkReqWrRmt_41 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[42]) begin
                    cntLkReqWrRmt_42 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[43]) begin
                    cntLkReqWrRmt_43 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[44]) begin
                    cntLkReqWrRmt_44 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[45]) begin
                    cntLkReqWrRmt_45 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[46]) begin
                    cntLkReqWrRmt_46 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[47]) begin
                    cntLkReqWrRmt_47 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[48]) begin
                    cntLkReqWrRmt_48 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[49]) begin
                    cntLkReqWrRmt_49 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[50]) begin
                    cntLkReqWrRmt_50 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[51]) begin
                    cntLkReqWrRmt_51 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[52]) begin
                    cntLkReqWrRmt_52 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[53]) begin
                    cntLkReqWrRmt_53 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[54]) begin
                    cntLkReqWrRmt_54 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[55]) begin
                    cntLkReqWrRmt_55 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[56]) begin
                    cntLkReqWrRmt_56 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[57]) begin
                    cntLkReqWrRmt_57 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[58]) begin
                    cntLkReqWrRmt_58 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[59]) begin
                    cntLkReqWrRmt_59 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[60]) begin
                    cntLkReqWrRmt_60 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[61]) begin
                    cntLkReqWrRmt_61 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[62]) begin
                    cntLkReqWrRmt_62 <= _zz_cntLkReqWrRmt_0_1;
                  end
                  if(_zz_85[63]) begin
                    cntLkReqWrRmt_63 <= _zz_cntLkReqWrRmt_0_1;
                  end
                end
              endcase
            end
          end
          if(when_TxnManCS_l128) begin
            if(_zz_86[0]) begin
              rReqDone_0 <= 1'b1;
            end
            if(_zz_86[1]) begin
              rReqDone_1 <= 1'b1;
            end
            if(_zz_86[2]) begin
              rReqDone_2 <= 1'b1;
            end
            if(_zz_86[3]) begin
              rReqDone_3 <= 1'b1;
            end
            if(_zz_86[4]) begin
              rReqDone_4 <= 1'b1;
            end
            if(_zz_86[5]) begin
              rReqDone_5 <= 1'b1;
            end
            if(_zz_86[6]) begin
              rReqDone_6 <= 1'b1;
            end
            if(_zz_86[7]) begin
              rReqDone_7 <= 1'b1;
            end
            if(_zz_86[8]) begin
              rReqDone_8 <= 1'b1;
            end
            if(_zz_86[9]) begin
              rReqDone_9 <= 1'b1;
            end
            if(_zz_86[10]) begin
              rReqDone_10 <= 1'b1;
            end
            if(_zz_86[11]) begin
              rReqDone_11 <= 1'b1;
            end
            if(_zz_86[12]) begin
              rReqDone_12 <= 1'b1;
            end
            if(_zz_86[13]) begin
              rReqDone_13 <= 1'b1;
            end
            if(_zz_86[14]) begin
              rReqDone_14 <= 1'b1;
            end
            if(_zz_86[15]) begin
              rReqDone_15 <= 1'b1;
            end
            if(_zz_86[16]) begin
              rReqDone_16 <= 1'b1;
            end
            if(_zz_86[17]) begin
              rReqDone_17 <= 1'b1;
            end
            if(_zz_86[18]) begin
              rReqDone_18 <= 1'b1;
            end
            if(_zz_86[19]) begin
              rReqDone_19 <= 1'b1;
            end
            if(_zz_86[20]) begin
              rReqDone_20 <= 1'b1;
            end
            if(_zz_86[21]) begin
              rReqDone_21 <= 1'b1;
            end
            if(_zz_86[22]) begin
              rReqDone_22 <= 1'b1;
            end
            if(_zz_86[23]) begin
              rReqDone_23 <= 1'b1;
            end
            if(_zz_86[24]) begin
              rReqDone_24 <= 1'b1;
            end
            if(_zz_86[25]) begin
              rReqDone_25 <= 1'b1;
            end
            if(_zz_86[26]) begin
              rReqDone_26 <= 1'b1;
            end
            if(_zz_86[27]) begin
              rReqDone_27 <= 1'b1;
            end
            if(_zz_86[28]) begin
              rReqDone_28 <= 1'b1;
            end
            if(_zz_86[29]) begin
              rReqDone_29 <= 1'b1;
            end
            if(_zz_86[30]) begin
              rReqDone_30 <= 1'b1;
            end
            if(_zz_86[31]) begin
              rReqDone_31 <= 1'b1;
            end
            if(_zz_86[32]) begin
              rReqDone_32 <= 1'b1;
            end
            if(_zz_86[33]) begin
              rReqDone_33 <= 1'b1;
            end
            if(_zz_86[34]) begin
              rReqDone_34 <= 1'b1;
            end
            if(_zz_86[35]) begin
              rReqDone_35 <= 1'b1;
            end
            if(_zz_86[36]) begin
              rReqDone_36 <= 1'b1;
            end
            if(_zz_86[37]) begin
              rReqDone_37 <= 1'b1;
            end
            if(_zz_86[38]) begin
              rReqDone_38 <= 1'b1;
            end
            if(_zz_86[39]) begin
              rReqDone_39 <= 1'b1;
            end
            if(_zz_86[40]) begin
              rReqDone_40 <= 1'b1;
            end
            if(_zz_86[41]) begin
              rReqDone_41 <= 1'b1;
            end
            if(_zz_86[42]) begin
              rReqDone_42 <= 1'b1;
            end
            if(_zz_86[43]) begin
              rReqDone_43 <= 1'b1;
            end
            if(_zz_86[44]) begin
              rReqDone_44 <= 1'b1;
            end
            if(_zz_86[45]) begin
              rReqDone_45 <= 1'b1;
            end
            if(_zz_86[46]) begin
              rReqDone_46 <= 1'b1;
            end
            if(_zz_86[47]) begin
              rReqDone_47 <= 1'b1;
            end
            if(_zz_86[48]) begin
              rReqDone_48 <= 1'b1;
            end
            if(_zz_86[49]) begin
              rReqDone_49 <= 1'b1;
            end
            if(_zz_86[50]) begin
              rReqDone_50 <= 1'b1;
            end
            if(_zz_86[51]) begin
              rReqDone_51 <= 1'b1;
            end
            if(_zz_86[52]) begin
              rReqDone_52 <= 1'b1;
            end
            if(_zz_86[53]) begin
              rReqDone_53 <= 1'b1;
            end
            if(_zz_86[54]) begin
              rReqDone_54 <= 1'b1;
            end
            if(_zz_86[55]) begin
              rReqDone_55 <= 1'b1;
            end
            if(_zz_86[56]) begin
              rReqDone_56 <= 1'b1;
            end
            if(_zz_86[57]) begin
              rReqDone_57 <= 1'b1;
            end
            if(_zz_86[58]) begin
              rReqDone_58 <= 1'b1;
            end
            if(_zz_86[59]) begin
              rReqDone_59 <= 1'b1;
            end
            if(_zz_86[60]) begin
              rReqDone_60 <= 1'b1;
            end
            if(_zz_86[61]) begin
              rReqDone_61 <= 1'b1;
            end
            if(_zz_86[62]) begin
              rReqDone_62 <= 1'b1;
            end
            if(_zz_86[63]) begin
              rReqDone_63 <= 1'b1;
            end
            compLkReq_reqIdx <= 6'h0;
          end
        end
        default : begin
        end
      endcase
      compLkRespLoc_stateReg <= compLkRespLoc_stateNext;
      case(compLkRespLoc_stateReg)
        compLkRespLoc_enumDef_WAIT_RESP : begin
          if(io_lkRespLoc_fire_3) begin
            case(io_lkRespLoc_payload_respType)
              LockRespType_grant : begin
                if(_zz_88) begin
                  cntLkRespLoc_0 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_89) begin
                  cntLkRespLoc_1 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_90) begin
                  cntLkRespLoc_2 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_91) begin
                  cntLkRespLoc_3 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_92) begin
                  cntLkRespLoc_4 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_93) begin
                  cntLkRespLoc_5 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_94) begin
                  cntLkRespLoc_6 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_95) begin
                  cntLkRespLoc_7 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_96) begin
                  cntLkRespLoc_8 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_97) begin
                  cntLkRespLoc_9 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_98) begin
                  cntLkRespLoc_10 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_99) begin
                  cntLkRespLoc_11 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_100) begin
                  cntLkRespLoc_12 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_101) begin
                  cntLkRespLoc_13 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_102) begin
                  cntLkRespLoc_14 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_103) begin
                  cntLkRespLoc_15 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_104) begin
                  cntLkRespLoc_16 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_105) begin
                  cntLkRespLoc_17 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_106) begin
                  cntLkRespLoc_18 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_107) begin
                  cntLkRespLoc_19 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_108) begin
                  cntLkRespLoc_20 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_109) begin
                  cntLkRespLoc_21 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_110) begin
                  cntLkRespLoc_22 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_111) begin
                  cntLkRespLoc_23 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_112) begin
                  cntLkRespLoc_24 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_113) begin
                  cntLkRespLoc_25 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_114) begin
                  cntLkRespLoc_26 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_115) begin
                  cntLkRespLoc_27 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_116) begin
                  cntLkRespLoc_28 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_117) begin
                  cntLkRespLoc_29 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_118) begin
                  cntLkRespLoc_30 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_119) begin
                  cntLkRespLoc_31 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_120) begin
                  cntLkRespLoc_32 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_121) begin
                  cntLkRespLoc_33 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_122) begin
                  cntLkRespLoc_34 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_123) begin
                  cntLkRespLoc_35 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_124) begin
                  cntLkRespLoc_36 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_125) begin
                  cntLkRespLoc_37 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_126) begin
                  cntLkRespLoc_38 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_127) begin
                  cntLkRespLoc_39 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_128) begin
                  cntLkRespLoc_40 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_129) begin
                  cntLkRespLoc_41 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_130) begin
                  cntLkRespLoc_42 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_131) begin
                  cntLkRespLoc_43 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_132) begin
                  cntLkRespLoc_44 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_133) begin
                  cntLkRespLoc_45 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_134) begin
                  cntLkRespLoc_46 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_135) begin
                  cntLkRespLoc_47 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_136) begin
                  cntLkRespLoc_48 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_137) begin
                  cntLkRespLoc_49 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_138) begin
                  cntLkRespLoc_50 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_139) begin
                  cntLkRespLoc_51 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_140) begin
                  cntLkRespLoc_52 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_141) begin
                  cntLkRespLoc_53 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_142) begin
                  cntLkRespLoc_54 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_143) begin
                  cntLkRespLoc_55 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_144) begin
                  cntLkRespLoc_56 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_145) begin
                  cntLkRespLoc_57 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_146) begin
                  cntLkRespLoc_58 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_147) begin
                  cntLkRespLoc_59 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_148) begin
                  cntLkRespLoc_60 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_149) begin
                  cntLkRespLoc_61 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_150) begin
                  cntLkRespLoc_62 <= _zz_cntLkRespLoc_0_1;
                end
                if(_zz_151) begin
                  cntLkRespLoc_63 <= _zz_cntLkRespLoc_0_1;
                end
                if(when_TxnManCS_l179) begin
                  if(_zz_6[0]) begin
                    cntLkHoldLoc_0 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[1]) begin
                    cntLkHoldLoc_1 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[2]) begin
                    cntLkHoldLoc_2 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[3]) begin
                    cntLkHoldLoc_3 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[4]) begin
                    cntLkHoldLoc_4 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[5]) begin
                    cntLkHoldLoc_5 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[6]) begin
                    cntLkHoldLoc_6 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[7]) begin
                    cntLkHoldLoc_7 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[8]) begin
                    cntLkHoldLoc_8 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[9]) begin
                    cntLkHoldLoc_9 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[10]) begin
                    cntLkHoldLoc_10 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[11]) begin
                    cntLkHoldLoc_11 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[12]) begin
                    cntLkHoldLoc_12 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[13]) begin
                    cntLkHoldLoc_13 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[14]) begin
                    cntLkHoldLoc_14 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[15]) begin
                    cntLkHoldLoc_15 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[16]) begin
                    cntLkHoldLoc_16 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[17]) begin
                    cntLkHoldLoc_17 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[18]) begin
                    cntLkHoldLoc_18 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[19]) begin
                    cntLkHoldLoc_19 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[20]) begin
                    cntLkHoldLoc_20 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[21]) begin
                    cntLkHoldLoc_21 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[22]) begin
                    cntLkHoldLoc_22 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[23]) begin
                    cntLkHoldLoc_23 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[24]) begin
                    cntLkHoldLoc_24 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[25]) begin
                    cntLkHoldLoc_25 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[26]) begin
                    cntLkHoldLoc_26 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[27]) begin
                    cntLkHoldLoc_27 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[28]) begin
                    cntLkHoldLoc_28 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[29]) begin
                    cntLkHoldLoc_29 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[30]) begin
                    cntLkHoldLoc_30 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[31]) begin
                    cntLkHoldLoc_31 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[32]) begin
                    cntLkHoldLoc_32 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[33]) begin
                    cntLkHoldLoc_33 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[34]) begin
                    cntLkHoldLoc_34 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[35]) begin
                    cntLkHoldLoc_35 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[36]) begin
                    cntLkHoldLoc_36 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[37]) begin
                    cntLkHoldLoc_37 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[38]) begin
                    cntLkHoldLoc_38 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[39]) begin
                    cntLkHoldLoc_39 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[40]) begin
                    cntLkHoldLoc_40 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[41]) begin
                    cntLkHoldLoc_41 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[42]) begin
                    cntLkHoldLoc_42 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[43]) begin
                    cntLkHoldLoc_43 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[44]) begin
                    cntLkHoldLoc_44 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[45]) begin
                    cntLkHoldLoc_45 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[46]) begin
                    cntLkHoldLoc_46 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[47]) begin
                    cntLkHoldLoc_47 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[48]) begin
                    cntLkHoldLoc_48 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[49]) begin
                    cntLkHoldLoc_49 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[50]) begin
                    cntLkHoldLoc_50 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[51]) begin
                    cntLkHoldLoc_51 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[52]) begin
                    cntLkHoldLoc_52 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[53]) begin
                    cntLkHoldLoc_53 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[54]) begin
                    cntLkHoldLoc_54 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[55]) begin
                    cntLkHoldLoc_55 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[56]) begin
                    cntLkHoldLoc_56 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[57]) begin
                    cntLkHoldLoc_57 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[58]) begin
                    cntLkHoldLoc_58 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[59]) begin
                    cntLkHoldLoc_59 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[60]) begin
                    cntLkHoldLoc_60 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[61]) begin
                    cntLkHoldLoc_61 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[62]) begin
                    cntLkHoldLoc_62 <= _zz_cntLkHoldLoc_0_1;
                  end
                  if(_zz_6[63]) begin
                    cntLkHoldLoc_63 <= _zz_cntLkHoldLoc_0_1;
                  end
                end
                case(io_lkRespLoc_payload_lkType)
                  LkT_rd : begin
                  end
                  LkT_wr : begin
                    if(_zz_153) begin
                      cntLkHoldWrLoc_0 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_154) begin
                      cntLkHoldWrLoc_1 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_155) begin
                      cntLkHoldWrLoc_2 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_156) begin
                      cntLkHoldWrLoc_3 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_157) begin
                      cntLkHoldWrLoc_4 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_158) begin
                      cntLkHoldWrLoc_5 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_159) begin
                      cntLkHoldWrLoc_6 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_160) begin
                      cntLkHoldWrLoc_7 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_161) begin
                      cntLkHoldWrLoc_8 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_162) begin
                      cntLkHoldWrLoc_9 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_163) begin
                      cntLkHoldWrLoc_10 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_164) begin
                      cntLkHoldWrLoc_11 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_165) begin
                      cntLkHoldWrLoc_12 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_166) begin
                      cntLkHoldWrLoc_13 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_167) begin
                      cntLkHoldWrLoc_14 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_168) begin
                      cntLkHoldWrLoc_15 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_169) begin
                      cntLkHoldWrLoc_16 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_170) begin
                      cntLkHoldWrLoc_17 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_171) begin
                      cntLkHoldWrLoc_18 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_172) begin
                      cntLkHoldWrLoc_19 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_173) begin
                      cntLkHoldWrLoc_20 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_174) begin
                      cntLkHoldWrLoc_21 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_175) begin
                      cntLkHoldWrLoc_22 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_176) begin
                      cntLkHoldWrLoc_23 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_177) begin
                      cntLkHoldWrLoc_24 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_178) begin
                      cntLkHoldWrLoc_25 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_179) begin
                      cntLkHoldWrLoc_26 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_180) begin
                      cntLkHoldWrLoc_27 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_181) begin
                      cntLkHoldWrLoc_28 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_182) begin
                      cntLkHoldWrLoc_29 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_183) begin
                      cntLkHoldWrLoc_30 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_184) begin
                      cntLkHoldWrLoc_31 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_185) begin
                      cntLkHoldWrLoc_32 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_186) begin
                      cntLkHoldWrLoc_33 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_187) begin
                      cntLkHoldWrLoc_34 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_188) begin
                      cntLkHoldWrLoc_35 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_189) begin
                      cntLkHoldWrLoc_36 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_190) begin
                      cntLkHoldWrLoc_37 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_191) begin
                      cntLkHoldWrLoc_38 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_192) begin
                      cntLkHoldWrLoc_39 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_193) begin
                      cntLkHoldWrLoc_40 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_194) begin
                      cntLkHoldWrLoc_41 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_195) begin
                      cntLkHoldWrLoc_42 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_196) begin
                      cntLkHoldWrLoc_43 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_197) begin
                      cntLkHoldWrLoc_44 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_198) begin
                      cntLkHoldWrLoc_45 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_199) begin
                      cntLkHoldWrLoc_46 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_200) begin
                      cntLkHoldWrLoc_47 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_201) begin
                      cntLkHoldWrLoc_48 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_202) begin
                      cntLkHoldWrLoc_49 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_203) begin
                      cntLkHoldWrLoc_50 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_204) begin
                      cntLkHoldWrLoc_51 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_205) begin
                      cntLkHoldWrLoc_52 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_206) begin
                      cntLkHoldWrLoc_53 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_207) begin
                      cntLkHoldWrLoc_54 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_208) begin
                      cntLkHoldWrLoc_55 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_209) begin
                      cntLkHoldWrLoc_56 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_210) begin
                      cntLkHoldWrLoc_57 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_211) begin
                      cntLkHoldWrLoc_58 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_212) begin
                      cntLkHoldWrLoc_59 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_213) begin
                      cntLkHoldWrLoc_60 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_214) begin
                      cntLkHoldWrLoc_61 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_215) begin
                      cntLkHoldWrLoc_62 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                    if(_zz_216) begin
                      cntLkHoldWrLoc_63 <= _zz_cntLkHoldWrLoc_0_1;
                    end
                  end
                  LkT_raw : begin
                    if(_zz_153) begin
                      cntLkHoldWrLoc_0 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_154) begin
                      cntLkHoldWrLoc_1 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_155) begin
                      cntLkHoldWrLoc_2 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_156) begin
                      cntLkHoldWrLoc_3 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_157) begin
                      cntLkHoldWrLoc_4 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_158) begin
                      cntLkHoldWrLoc_5 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_159) begin
                      cntLkHoldWrLoc_6 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_160) begin
                      cntLkHoldWrLoc_7 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_161) begin
                      cntLkHoldWrLoc_8 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_162) begin
                      cntLkHoldWrLoc_9 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_163) begin
                      cntLkHoldWrLoc_10 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_164) begin
                      cntLkHoldWrLoc_11 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_165) begin
                      cntLkHoldWrLoc_12 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_166) begin
                      cntLkHoldWrLoc_13 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_167) begin
                      cntLkHoldWrLoc_14 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_168) begin
                      cntLkHoldWrLoc_15 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_169) begin
                      cntLkHoldWrLoc_16 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_170) begin
                      cntLkHoldWrLoc_17 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_171) begin
                      cntLkHoldWrLoc_18 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_172) begin
                      cntLkHoldWrLoc_19 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_173) begin
                      cntLkHoldWrLoc_20 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_174) begin
                      cntLkHoldWrLoc_21 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_175) begin
                      cntLkHoldWrLoc_22 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_176) begin
                      cntLkHoldWrLoc_23 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_177) begin
                      cntLkHoldWrLoc_24 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_178) begin
                      cntLkHoldWrLoc_25 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_179) begin
                      cntLkHoldWrLoc_26 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_180) begin
                      cntLkHoldWrLoc_27 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_181) begin
                      cntLkHoldWrLoc_28 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_182) begin
                      cntLkHoldWrLoc_29 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_183) begin
                      cntLkHoldWrLoc_30 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_184) begin
                      cntLkHoldWrLoc_31 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_185) begin
                      cntLkHoldWrLoc_32 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_186) begin
                      cntLkHoldWrLoc_33 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_187) begin
                      cntLkHoldWrLoc_34 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_188) begin
                      cntLkHoldWrLoc_35 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_189) begin
                      cntLkHoldWrLoc_36 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_190) begin
                      cntLkHoldWrLoc_37 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_191) begin
                      cntLkHoldWrLoc_38 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_192) begin
                      cntLkHoldWrLoc_39 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_193) begin
                      cntLkHoldWrLoc_40 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_194) begin
                      cntLkHoldWrLoc_41 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_195) begin
                      cntLkHoldWrLoc_42 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_196) begin
                      cntLkHoldWrLoc_43 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_197) begin
                      cntLkHoldWrLoc_44 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_198) begin
                      cntLkHoldWrLoc_45 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_199) begin
                      cntLkHoldWrLoc_46 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_200) begin
                      cntLkHoldWrLoc_47 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_201) begin
                      cntLkHoldWrLoc_48 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_202) begin
                      cntLkHoldWrLoc_49 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_203) begin
                      cntLkHoldWrLoc_50 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_204) begin
                      cntLkHoldWrLoc_51 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_205) begin
                      cntLkHoldWrLoc_52 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_206) begin
                      cntLkHoldWrLoc_53 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_207) begin
                      cntLkHoldWrLoc_54 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_208) begin
                      cntLkHoldWrLoc_55 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_209) begin
                      cntLkHoldWrLoc_56 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_210) begin
                      cntLkHoldWrLoc_57 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_211) begin
                      cntLkHoldWrLoc_58 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_212) begin
                      cntLkHoldWrLoc_59 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_213) begin
                      cntLkHoldWrLoc_60 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_214) begin
                      cntLkHoldWrLoc_61 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_215) begin
                      cntLkHoldWrLoc_62 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                    if(_zz_216) begin
                      cntLkHoldWrLoc_63 <= _zz_cntLkHoldWrLoc_0_2;
                    end
                  end
                  default : begin
                  end
                endcase
              end
              LockRespType_waiting : begin
                if(_zz_7[0]) begin
                  cntLkWaitLoc_0 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[1]) begin
                  cntLkWaitLoc_1 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[2]) begin
                  cntLkWaitLoc_2 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[3]) begin
                  cntLkWaitLoc_3 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[4]) begin
                  cntLkWaitLoc_4 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[5]) begin
                  cntLkWaitLoc_5 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[6]) begin
                  cntLkWaitLoc_6 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[7]) begin
                  cntLkWaitLoc_7 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[8]) begin
                  cntLkWaitLoc_8 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[9]) begin
                  cntLkWaitLoc_9 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[10]) begin
                  cntLkWaitLoc_10 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[11]) begin
                  cntLkWaitLoc_11 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[12]) begin
                  cntLkWaitLoc_12 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[13]) begin
                  cntLkWaitLoc_13 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[14]) begin
                  cntLkWaitLoc_14 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[15]) begin
                  cntLkWaitLoc_15 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[16]) begin
                  cntLkWaitLoc_16 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[17]) begin
                  cntLkWaitLoc_17 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[18]) begin
                  cntLkWaitLoc_18 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[19]) begin
                  cntLkWaitLoc_19 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[20]) begin
                  cntLkWaitLoc_20 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[21]) begin
                  cntLkWaitLoc_21 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[22]) begin
                  cntLkWaitLoc_22 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[23]) begin
                  cntLkWaitLoc_23 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[24]) begin
                  cntLkWaitLoc_24 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[25]) begin
                  cntLkWaitLoc_25 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[26]) begin
                  cntLkWaitLoc_26 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[27]) begin
                  cntLkWaitLoc_27 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[28]) begin
                  cntLkWaitLoc_28 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[29]) begin
                  cntLkWaitLoc_29 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[30]) begin
                  cntLkWaitLoc_30 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[31]) begin
                  cntLkWaitLoc_31 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[32]) begin
                  cntLkWaitLoc_32 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[33]) begin
                  cntLkWaitLoc_33 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[34]) begin
                  cntLkWaitLoc_34 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[35]) begin
                  cntLkWaitLoc_35 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[36]) begin
                  cntLkWaitLoc_36 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[37]) begin
                  cntLkWaitLoc_37 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[38]) begin
                  cntLkWaitLoc_38 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[39]) begin
                  cntLkWaitLoc_39 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[40]) begin
                  cntLkWaitLoc_40 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[41]) begin
                  cntLkWaitLoc_41 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[42]) begin
                  cntLkWaitLoc_42 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[43]) begin
                  cntLkWaitLoc_43 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[44]) begin
                  cntLkWaitLoc_44 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[45]) begin
                  cntLkWaitLoc_45 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[46]) begin
                  cntLkWaitLoc_46 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[47]) begin
                  cntLkWaitLoc_47 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[48]) begin
                  cntLkWaitLoc_48 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[49]) begin
                  cntLkWaitLoc_49 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[50]) begin
                  cntLkWaitLoc_50 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[51]) begin
                  cntLkWaitLoc_51 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[52]) begin
                  cntLkWaitLoc_52 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[53]) begin
                  cntLkWaitLoc_53 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[54]) begin
                  cntLkWaitLoc_54 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[55]) begin
                  cntLkWaitLoc_55 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[56]) begin
                  cntLkWaitLoc_56 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[57]) begin
                  cntLkWaitLoc_57 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[58]) begin
                  cntLkWaitLoc_58 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[59]) begin
                  cntLkWaitLoc_59 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[60]) begin
                  cntLkWaitLoc_60 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[61]) begin
                  cntLkWaitLoc_61 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[62]) begin
                  cntLkWaitLoc_62 <= _zz_cntLkWaitLoc_0_1;
                end
                if(_zz_7[63]) begin
                  cntLkWaitLoc_63 <= _zz_cntLkWaitLoc_0_1;
                end
              end
              LockRespType_abort : begin
                if(_zz_217[0]) begin
                  rAbort_0 <= 1'b1;
                end
                if(_zz_217[1]) begin
                  rAbort_1 <= 1'b1;
                end
                if(_zz_217[2]) begin
                  rAbort_2 <= 1'b1;
                end
                if(_zz_217[3]) begin
                  rAbort_3 <= 1'b1;
                end
                if(_zz_217[4]) begin
                  rAbort_4 <= 1'b1;
                end
                if(_zz_217[5]) begin
                  rAbort_5 <= 1'b1;
                end
                if(_zz_217[6]) begin
                  rAbort_6 <= 1'b1;
                end
                if(_zz_217[7]) begin
                  rAbort_7 <= 1'b1;
                end
                if(_zz_217[8]) begin
                  rAbort_8 <= 1'b1;
                end
                if(_zz_217[9]) begin
                  rAbort_9 <= 1'b1;
                end
                if(_zz_217[10]) begin
                  rAbort_10 <= 1'b1;
                end
                if(_zz_217[11]) begin
                  rAbort_11 <= 1'b1;
                end
                if(_zz_217[12]) begin
                  rAbort_12 <= 1'b1;
                end
                if(_zz_217[13]) begin
                  rAbort_13 <= 1'b1;
                end
                if(_zz_217[14]) begin
                  rAbort_14 <= 1'b1;
                end
                if(_zz_217[15]) begin
                  rAbort_15 <= 1'b1;
                end
                if(_zz_217[16]) begin
                  rAbort_16 <= 1'b1;
                end
                if(_zz_217[17]) begin
                  rAbort_17 <= 1'b1;
                end
                if(_zz_217[18]) begin
                  rAbort_18 <= 1'b1;
                end
                if(_zz_217[19]) begin
                  rAbort_19 <= 1'b1;
                end
                if(_zz_217[20]) begin
                  rAbort_20 <= 1'b1;
                end
                if(_zz_217[21]) begin
                  rAbort_21 <= 1'b1;
                end
                if(_zz_217[22]) begin
                  rAbort_22 <= 1'b1;
                end
                if(_zz_217[23]) begin
                  rAbort_23 <= 1'b1;
                end
                if(_zz_217[24]) begin
                  rAbort_24 <= 1'b1;
                end
                if(_zz_217[25]) begin
                  rAbort_25 <= 1'b1;
                end
                if(_zz_217[26]) begin
                  rAbort_26 <= 1'b1;
                end
                if(_zz_217[27]) begin
                  rAbort_27 <= 1'b1;
                end
                if(_zz_217[28]) begin
                  rAbort_28 <= 1'b1;
                end
                if(_zz_217[29]) begin
                  rAbort_29 <= 1'b1;
                end
                if(_zz_217[30]) begin
                  rAbort_30 <= 1'b1;
                end
                if(_zz_217[31]) begin
                  rAbort_31 <= 1'b1;
                end
                if(_zz_217[32]) begin
                  rAbort_32 <= 1'b1;
                end
                if(_zz_217[33]) begin
                  rAbort_33 <= 1'b1;
                end
                if(_zz_217[34]) begin
                  rAbort_34 <= 1'b1;
                end
                if(_zz_217[35]) begin
                  rAbort_35 <= 1'b1;
                end
                if(_zz_217[36]) begin
                  rAbort_36 <= 1'b1;
                end
                if(_zz_217[37]) begin
                  rAbort_37 <= 1'b1;
                end
                if(_zz_217[38]) begin
                  rAbort_38 <= 1'b1;
                end
                if(_zz_217[39]) begin
                  rAbort_39 <= 1'b1;
                end
                if(_zz_217[40]) begin
                  rAbort_40 <= 1'b1;
                end
                if(_zz_217[41]) begin
                  rAbort_41 <= 1'b1;
                end
                if(_zz_217[42]) begin
                  rAbort_42 <= 1'b1;
                end
                if(_zz_217[43]) begin
                  rAbort_43 <= 1'b1;
                end
                if(_zz_217[44]) begin
                  rAbort_44 <= 1'b1;
                end
                if(_zz_217[45]) begin
                  rAbort_45 <= 1'b1;
                end
                if(_zz_217[46]) begin
                  rAbort_46 <= 1'b1;
                end
                if(_zz_217[47]) begin
                  rAbort_47 <= 1'b1;
                end
                if(_zz_217[48]) begin
                  rAbort_48 <= 1'b1;
                end
                if(_zz_217[49]) begin
                  rAbort_49 <= 1'b1;
                end
                if(_zz_217[50]) begin
                  rAbort_50 <= 1'b1;
                end
                if(_zz_217[51]) begin
                  rAbort_51 <= 1'b1;
                end
                if(_zz_217[52]) begin
                  rAbort_52 <= 1'b1;
                end
                if(_zz_217[53]) begin
                  rAbort_53 <= 1'b1;
                end
                if(_zz_217[54]) begin
                  rAbort_54 <= 1'b1;
                end
                if(_zz_217[55]) begin
                  rAbort_55 <= 1'b1;
                end
                if(_zz_217[56]) begin
                  rAbort_56 <= 1'b1;
                end
                if(_zz_217[57]) begin
                  rAbort_57 <= 1'b1;
                end
                if(_zz_217[58]) begin
                  rAbort_58 <= 1'b1;
                end
                if(_zz_217[59]) begin
                  rAbort_59 <= 1'b1;
                end
                if(_zz_217[60]) begin
                  rAbort_60 <= 1'b1;
                end
                if(_zz_217[61]) begin
                  rAbort_61 <= 1'b1;
                end
                if(_zz_217[62]) begin
                  rAbort_62 <= 1'b1;
                end
                if(_zz_217[63]) begin
                  rAbort_63 <= 1'b1;
                end
                if(_zz_88) begin
                  cntLkRespLoc_0 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_89) begin
                  cntLkRespLoc_1 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_90) begin
                  cntLkRespLoc_2 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_91) begin
                  cntLkRespLoc_3 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_92) begin
                  cntLkRespLoc_4 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_93) begin
                  cntLkRespLoc_5 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_94) begin
                  cntLkRespLoc_6 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_95) begin
                  cntLkRespLoc_7 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_96) begin
                  cntLkRespLoc_8 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_97) begin
                  cntLkRespLoc_9 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_98) begin
                  cntLkRespLoc_10 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_99) begin
                  cntLkRespLoc_11 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_100) begin
                  cntLkRespLoc_12 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_101) begin
                  cntLkRespLoc_13 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_102) begin
                  cntLkRespLoc_14 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_103) begin
                  cntLkRespLoc_15 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_104) begin
                  cntLkRespLoc_16 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_105) begin
                  cntLkRespLoc_17 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_106) begin
                  cntLkRespLoc_18 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_107) begin
                  cntLkRespLoc_19 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_108) begin
                  cntLkRespLoc_20 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_109) begin
                  cntLkRespLoc_21 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_110) begin
                  cntLkRespLoc_22 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_111) begin
                  cntLkRespLoc_23 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_112) begin
                  cntLkRespLoc_24 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_113) begin
                  cntLkRespLoc_25 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_114) begin
                  cntLkRespLoc_26 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_115) begin
                  cntLkRespLoc_27 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_116) begin
                  cntLkRespLoc_28 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_117) begin
                  cntLkRespLoc_29 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_118) begin
                  cntLkRespLoc_30 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_119) begin
                  cntLkRespLoc_31 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_120) begin
                  cntLkRespLoc_32 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_121) begin
                  cntLkRespLoc_33 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_122) begin
                  cntLkRespLoc_34 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_123) begin
                  cntLkRespLoc_35 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_124) begin
                  cntLkRespLoc_36 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_125) begin
                  cntLkRespLoc_37 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_126) begin
                  cntLkRespLoc_38 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_127) begin
                  cntLkRespLoc_39 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_128) begin
                  cntLkRespLoc_40 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_129) begin
                  cntLkRespLoc_41 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_130) begin
                  cntLkRespLoc_42 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_131) begin
                  cntLkRespLoc_43 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_132) begin
                  cntLkRespLoc_44 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_133) begin
                  cntLkRespLoc_45 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_134) begin
                  cntLkRespLoc_46 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_135) begin
                  cntLkRespLoc_47 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_136) begin
                  cntLkRespLoc_48 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_137) begin
                  cntLkRespLoc_49 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_138) begin
                  cntLkRespLoc_50 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_139) begin
                  cntLkRespLoc_51 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_140) begin
                  cntLkRespLoc_52 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_141) begin
                  cntLkRespLoc_53 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_142) begin
                  cntLkRespLoc_54 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_143) begin
                  cntLkRespLoc_55 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_144) begin
                  cntLkRespLoc_56 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_145) begin
                  cntLkRespLoc_57 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_146) begin
                  cntLkRespLoc_58 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_147) begin
                  cntLkRespLoc_59 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_148) begin
                  cntLkRespLoc_60 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_149) begin
                  cntLkRespLoc_61 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_150) begin
                  cntLkRespLoc_62 <= _zz_cntLkRespLoc_0_2;
                end
                if(_zz_151) begin
                  cntLkRespLoc_63 <= _zz_cntLkRespLoc_0_2;
                end
                io_cntLockDenyLoc <= (io_cntLockDenyLoc + 32'h00000001);
              end
              default : begin
                if(_zz_5[0]) begin
                  cntRlseRespLoc_0 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[1]) begin
                  cntRlseRespLoc_1 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[2]) begin
                  cntRlseRespLoc_2 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[3]) begin
                  cntRlseRespLoc_3 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[4]) begin
                  cntRlseRespLoc_4 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[5]) begin
                  cntRlseRespLoc_5 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[6]) begin
                  cntRlseRespLoc_6 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[7]) begin
                  cntRlseRespLoc_7 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[8]) begin
                  cntRlseRespLoc_8 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[9]) begin
                  cntRlseRespLoc_9 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[10]) begin
                  cntRlseRespLoc_10 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[11]) begin
                  cntRlseRespLoc_11 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[12]) begin
                  cntRlseRespLoc_12 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[13]) begin
                  cntRlseRespLoc_13 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[14]) begin
                  cntRlseRespLoc_14 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[15]) begin
                  cntRlseRespLoc_15 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[16]) begin
                  cntRlseRespLoc_16 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[17]) begin
                  cntRlseRespLoc_17 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[18]) begin
                  cntRlseRespLoc_18 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[19]) begin
                  cntRlseRespLoc_19 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[20]) begin
                  cntRlseRespLoc_20 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[21]) begin
                  cntRlseRespLoc_21 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[22]) begin
                  cntRlseRespLoc_22 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[23]) begin
                  cntRlseRespLoc_23 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[24]) begin
                  cntRlseRespLoc_24 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[25]) begin
                  cntRlseRespLoc_25 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[26]) begin
                  cntRlseRespLoc_26 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[27]) begin
                  cntRlseRespLoc_27 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[28]) begin
                  cntRlseRespLoc_28 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[29]) begin
                  cntRlseRespLoc_29 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[30]) begin
                  cntRlseRespLoc_30 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[31]) begin
                  cntRlseRespLoc_31 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[32]) begin
                  cntRlseRespLoc_32 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[33]) begin
                  cntRlseRespLoc_33 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[34]) begin
                  cntRlseRespLoc_34 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[35]) begin
                  cntRlseRespLoc_35 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[36]) begin
                  cntRlseRespLoc_36 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[37]) begin
                  cntRlseRespLoc_37 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[38]) begin
                  cntRlseRespLoc_38 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[39]) begin
                  cntRlseRespLoc_39 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[40]) begin
                  cntRlseRespLoc_40 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[41]) begin
                  cntRlseRespLoc_41 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[42]) begin
                  cntRlseRespLoc_42 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[43]) begin
                  cntRlseRespLoc_43 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[44]) begin
                  cntRlseRespLoc_44 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[45]) begin
                  cntRlseRespLoc_45 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[46]) begin
                  cntRlseRespLoc_46 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[47]) begin
                  cntRlseRespLoc_47 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[48]) begin
                  cntRlseRespLoc_48 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[49]) begin
                  cntRlseRespLoc_49 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[50]) begin
                  cntRlseRespLoc_50 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[51]) begin
                  cntRlseRespLoc_51 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[52]) begin
                  cntRlseRespLoc_52 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[53]) begin
                  cntRlseRespLoc_53 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[54]) begin
                  cntRlseRespLoc_54 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[55]) begin
                  cntRlseRespLoc_55 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[56]) begin
                  cntRlseRespLoc_56 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[57]) begin
                  cntRlseRespLoc_57 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[58]) begin
                  cntRlseRespLoc_58 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[59]) begin
                  cntRlseRespLoc_59 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[60]) begin
                  cntRlseRespLoc_60 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[61]) begin
                  cntRlseRespLoc_61 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[62]) begin
                  cntRlseRespLoc_62 <= _zz_cntRlseRespLoc_0_1;
                end
                if(_zz_5[63]) begin
                  cntRlseRespLoc_63 <= _zz_cntRlseRespLoc_0_1;
                end
              end
            endcase
          end
        end
        compLkRespLoc_enumDef_LOCAL_RD_REQ : begin
        end
        default : begin
        end
      endcase
      compLkRespRmt_stateReg <= compLkRespRmt_stateNext;
      case(compLkRespRmt_stateReg)
        compLkRespRmt_enumDef_WAIT_RESP : begin
          if(io_lkRespRmt_fire_3) begin
            case(io_lkRespRmt_payload_respType)
              LockRespType_grant : begin
                if(_zz_219) begin
                  cntLkRespRmt_0 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_220) begin
                  cntLkRespRmt_1 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_221) begin
                  cntLkRespRmt_2 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_222) begin
                  cntLkRespRmt_3 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_223) begin
                  cntLkRespRmt_4 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_224) begin
                  cntLkRespRmt_5 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_225) begin
                  cntLkRespRmt_6 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_226) begin
                  cntLkRespRmt_7 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_227) begin
                  cntLkRespRmt_8 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_228) begin
                  cntLkRespRmt_9 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_229) begin
                  cntLkRespRmt_10 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_230) begin
                  cntLkRespRmt_11 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_231) begin
                  cntLkRespRmt_12 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_232) begin
                  cntLkRespRmt_13 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_233) begin
                  cntLkRespRmt_14 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_234) begin
                  cntLkRespRmt_15 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_235) begin
                  cntLkRespRmt_16 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_236) begin
                  cntLkRespRmt_17 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_237) begin
                  cntLkRespRmt_18 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_238) begin
                  cntLkRespRmt_19 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_239) begin
                  cntLkRespRmt_20 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_240) begin
                  cntLkRespRmt_21 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_241) begin
                  cntLkRespRmt_22 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_242) begin
                  cntLkRespRmt_23 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_243) begin
                  cntLkRespRmt_24 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_244) begin
                  cntLkRespRmt_25 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_245) begin
                  cntLkRespRmt_26 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_246) begin
                  cntLkRespRmt_27 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_247) begin
                  cntLkRespRmt_28 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_248) begin
                  cntLkRespRmt_29 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_249) begin
                  cntLkRespRmt_30 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_250) begin
                  cntLkRespRmt_31 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_251) begin
                  cntLkRespRmt_32 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_252) begin
                  cntLkRespRmt_33 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_253) begin
                  cntLkRespRmt_34 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_254) begin
                  cntLkRespRmt_35 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_255) begin
                  cntLkRespRmt_36 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_256) begin
                  cntLkRespRmt_37 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_257) begin
                  cntLkRespRmt_38 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_258) begin
                  cntLkRespRmt_39 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_259) begin
                  cntLkRespRmt_40 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_260) begin
                  cntLkRespRmt_41 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_261) begin
                  cntLkRespRmt_42 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_262) begin
                  cntLkRespRmt_43 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_263) begin
                  cntLkRespRmt_44 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_264) begin
                  cntLkRespRmt_45 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_265) begin
                  cntLkRespRmt_46 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_266) begin
                  cntLkRespRmt_47 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_267) begin
                  cntLkRespRmt_48 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_268) begin
                  cntLkRespRmt_49 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_269) begin
                  cntLkRespRmt_50 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_270) begin
                  cntLkRespRmt_51 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_271) begin
                  cntLkRespRmt_52 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_272) begin
                  cntLkRespRmt_53 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_273) begin
                  cntLkRespRmt_54 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_274) begin
                  cntLkRespRmt_55 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_275) begin
                  cntLkRespRmt_56 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_276) begin
                  cntLkRespRmt_57 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_277) begin
                  cntLkRespRmt_58 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_278) begin
                  cntLkRespRmt_59 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_279) begin
                  cntLkRespRmt_60 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_280) begin
                  cntLkRespRmt_61 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_281) begin
                  cntLkRespRmt_62 <= _zz_cntLkRespRmt_0_1;
                end
                if(_zz_282) begin
                  cntLkRespRmt_63 <= _zz_cntLkRespRmt_0_1;
                end
                if(when_TxnManCS_l272) begin
                  if(_zz_10[0]) begin
                    cntLkHoldRmt_0 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[1]) begin
                    cntLkHoldRmt_1 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[2]) begin
                    cntLkHoldRmt_2 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[3]) begin
                    cntLkHoldRmt_3 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[4]) begin
                    cntLkHoldRmt_4 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[5]) begin
                    cntLkHoldRmt_5 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[6]) begin
                    cntLkHoldRmt_6 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[7]) begin
                    cntLkHoldRmt_7 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[8]) begin
                    cntLkHoldRmt_8 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[9]) begin
                    cntLkHoldRmt_9 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[10]) begin
                    cntLkHoldRmt_10 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[11]) begin
                    cntLkHoldRmt_11 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[12]) begin
                    cntLkHoldRmt_12 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[13]) begin
                    cntLkHoldRmt_13 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[14]) begin
                    cntLkHoldRmt_14 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[15]) begin
                    cntLkHoldRmt_15 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[16]) begin
                    cntLkHoldRmt_16 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[17]) begin
                    cntLkHoldRmt_17 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[18]) begin
                    cntLkHoldRmt_18 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[19]) begin
                    cntLkHoldRmt_19 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[20]) begin
                    cntLkHoldRmt_20 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[21]) begin
                    cntLkHoldRmt_21 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[22]) begin
                    cntLkHoldRmt_22 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[23]) begin
                    cntLkHoldRmt_23 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[24]) begin
                    cntLkHoldRmt_24 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[25]) begin
                    cntLkHoldRmt_25 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[26]) begin
                    cntLkHoldRmt_26 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[27]) begin
                    cntLkHoldRmt_27 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[28]) begin
                    cntLkHoldRmt_28 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[29]) begin
                    cntLkHoldRmt_29 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[30]) begin
                    cntLkHoldRmt_30 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[31]) begin
                    cntLkHoldRmt_31 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[32]) begin
                    cntLkHoldRmt_32 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[33]) begin
                    cntLkHoldRmt_33 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[34]) begin
                    cntLkHoldRmt_34 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[35]) begin
                    cntLkHoldRmt_35 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[36]) begin
                    cntLkHoldRmt_36 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[37]) begin
                    cntLkHoldRmt_37 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[38]) begin
                    cntLkHoldRmt_38 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[39]) begin
                    cntLkHoldRmt_39 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[40]) begin
                    cntLkHoldRmt_40 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[41]) begin
                    cntLkHoldRmt_41 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[42]) begin
                    cntLkHoldRmt_42 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[43]) begin
                    cntLkHoldRmt_43 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[44]) begin
                    cntLkHoldRmt_44 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[45]) begin
                    cntLkHoldRmt_45 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[46]) begin
                    cntLkHoldRmt_46 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[47]) begin
                    cntLkHoldRmt_47 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[48]) begin
                    cntLkHoldRmt_48 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[49]) begin
                    cntLkHoldRmt_49 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[50]) begin
                    cntLkHoldRmt_50 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[51]) begin
                    cntLkHoldRmt_51 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[52]) begin
                    cntLkHoldRmt_52 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[53]) begin
                    cntLkHoldRmt_53 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[54]) begin
                    cntLkHoldRmt_54 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[55]) begin
                    cntLkHoldRmt_55 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[56]) begin
                    cntLkHoldRmt_56 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[57]) begin
                    cntLkHoldRmt_57 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[58]) begin
                    cntLkHoldRmt_58 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[59]) begin
                    cntLkHoldRmt_59 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[60]) begin
                    cntLkHoldRmt_60 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[61]) begin
                    cntLkHoldRmt_61 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[62]) begin
                    cntLkHoldRmt_62 <= _zz_cntLkHoldRmt_0_1;
                  end
                  if(_zz_10[63]) begin
                    cntLkHoldRmt_63 <= _zz_cntLkHoldRmt_0_1;
                  end
                end
                case(io_lkRespRmt_payload_lkType)
                  LkT_rd : begin
                  end
                  LkT_wr : begin
                    if(_zz_284) begin
                      cntLkHoldWrRmt_0 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_285) begin
                      cntLkHoldWrRmt_1 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_286) begin
                      cntLkHoldWrRmt_2 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_287) begin
                      cntLkHoldWrRmt_3 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_288) begin
                      cntLkHoldWrRmt_4 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_289) begin
                      cntLkHoldWrRmt_5 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_290) begin
                      cntLkHoldWrRmt_6 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_291) begin
                      cntLkHoldWrRmt_7 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_292) begin
                      cntLkHoldWrRmt_8 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_293) begin
                      cntLkHoldWrRmt_9 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_294) begin
                      cntLkHoldWrRmt_10 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_295) begin
                      cntLkHoldWrRmt_11 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_296) begin
                      cntLkHoldWrRmt_12 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_297) begin
                      cntLkHoldWrRmt_13 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_298) begin
                      cntLkHoldWrRmt_14 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_299) begin
                      cntLkHoldWrRmt_15 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_300) begin
                      cntLkHoldWrRmt_16 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_301) begin
                      cntLkHoldWrRmt_17 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_302) begin
                      cntLkHoldWrRmt_18 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_303) begin
                      cntLkHoldWrRmt_19 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_304) begin
                      cntLkHoldWrRmt_20 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_305) begin
                      cntLkHoldWrRmt_21 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_306) begin
                      cntLkHoldWrRmt_22 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_307) begin
                      cntLkHoldWrRmt_23 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_308) begin
                      cntLkHoldWrRmt_24 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_309) begin
                      cntLkHoldWrRmt_25 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_310) begin
                      cntLkHoldWrRmt_26 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_311) begin
                      cntLkHoldWrRmt_27 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_312) begin
                      cntLkHoldWrRmt_28 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_313) begin
                      cntLkHoldWrRmt_29 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_314) begin
                      cntLkHoldWrRmt_30 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_315) begin
                      cntLkHoldWrRmt_31 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_316) begin
                      cntLkHoldWrRmt_32 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_317) begin
                      cntLkHoldWrRmt_33 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_318) begin
                      cntLkHoldWrRmt_34 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_319) begin
                      cntLkHoldWrRmt_35 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_320) begin
                      cntLkHoldWrRmt_36 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_321) begin
                      cntLkHoldWrRmt_37 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_322) begin
                      cntLkHoldWrRmt_38 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_323) begin
                      cntLkHoldWrRmt_39 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_324) begin
                      cntLkHoldWrRmt_40 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_325) begin
                      cntLkHoldWrRmt_41 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_326) begin
                      cntLkHoldWrRmt_42 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_327) begin
                      cntLkHoldWrRmt_43 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_328) begin
                      cntLkHoldWrRmt_44 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_329) begin
                      cntLkHoldWrRmt_45 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_330) begin
                      cntLkHoldWrRmt_46 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_331) begin
                      cntLkHoldWrRmt_47 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_332) begin
                      cntLkHoldWrRmt_48 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_333) begin
                      cntLkHoldWrRmt_49 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_334) begin
                      cntLkHoldWrRmt_50 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_335) begin
                      cntLkHoldWrRmt_51 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_336) begin
                      cntLkHoldWrRmt_52 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_337) begin
                      cntLkHoldWrRmt_53 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_338) begin
                      cntLkHoldWrRmt_54 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_339) begin
                      cntLkHoldWrRmt_55 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_340) begin
                      cntLkHoldWrRmt_56 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_341) begin
                      cntLkHoldWrRmt_57 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_342) begin
                      cntLkHoldWrRmt_58 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_343) begin
                      cntLkHoldWrRmt_59 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_344) begin
                      cntLkHoldWrRmt_60 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_345) begin
                      cntLkHoldWrRmt_61 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_346) begin
                      cntLkHoldWrRmt_62 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                    if(_zz_347) begin
                      cntLkHoldWrRmt_63 <= _zz_cntLkHoldWrRmt_0_1;
                    end
                  end
                  LkT_raw : begin
                    if(_zz_284) begin
                      cntLkHoldWrRmt_0 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_285) begin
                      cntLkHoldWrRmt_1 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_286) begin
                      cntLkHoldWrRmt_2 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_287) begin
                      cntLkHoldWrRmt_3 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_288) begin
                      cntLkHoldWrRmt_4 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_289) begin
                      cntLkHoldWrRmt_5 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_290) begin
                      cntLkHoldWrRmt_6 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_291) begin
                      cntLkHoldWrRmt_7 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_292) begin
                      cntLkHoldWrRmt_8 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_293) begin
                      cntLkHoldWrRmt_9 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_294) begin
                      cntLkHoldWrRmt_10 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_295) begin
                      cntLkHoldWrRmt_11 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_296) begin
                      cntLkHoldWrRmt_12 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_297) begin
                      cntLkHoldWrRmt_13 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_298) begin
                      cntLkHoldWrRmt_14 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_299) begin
                      cntLkHoldWrRmt_15 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_300) begin
                      cntLkHoldWrRmt_16 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_301) begin
                      cntLkHoldWrRmt_17 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_302) begin
                      cntLkHoldWrRmt_18 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_303) begin
                      cntLkHoldWrRmt_19 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_304) begin
                      cntLkHoldWrRmt_20 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_305) begin
                      cntLkHoldWrRmt_21 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_306) begin
                      cntLkHoldWrRmt_22 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_307) begin
                      cntLkHoldWrRmt_23 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_308) begin
                      cntLkHoldWrRmt_24 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_309) begin
                      cntLkHoldWrRmt_25 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_310) begin
                      cntLkHoldWrRmt_26 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_311) begin
                      cntLkHoldWrRmt_27 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_312) begin
                      cntLkHoldWrRmt_28 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_313) begin
                      cntLkHoldWrRmt_29 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_314) begin
                      cntLkHoldWrRmt_30 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_315) begin
                      cntLkHoldWrRmt_31 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_316) begin
                      cntLkHoldWrRmt_32 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_317) begin
                      cntLkHoldWrRmt_33 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_318) begin
                      cntLkHoldWrRmt_34 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_319) begin
                      cntLkHoldWrRmt_35 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_320) begin
                      cntLkHoldWrRmt_36 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_321) begin
                      cntLkHoldWrRmt_37 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_322) begin
                      cntLkHoldWrRmt_38 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_323) begin
                      cntLkHoldWrRmt_39 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_324) begin
                      cntLkHoldWrRmt_40 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_325) begin
                      cntLkHoldWrRmt_41 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_326) begin
                      cntLkHoldWrRmt_42 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_327) begin
                      cntLkHoldWrRmt_43 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_328) begin
                      cntLkHoldWrRmt_44 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_329) begin
                      cntLkHoldWrRmt_45 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_330) begin
                      cntLkHoldWrRmt_46 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_331) begin
                      cntLkHoldWrRmt_47 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_332) begin
                      cntLkHoldWrRmt_48 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_333) begin
                      cntLkHoldWrRmt_49 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_334) begin
                      cntLkHoldWrRmt_50 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_335) begin
                      cntLkHoldWrRmt_51 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_336) begin
                      cntLkHoldWrRmt_52 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_337) begin
                      cntLkHoldWrRmt_53 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_338) begin
                      cntLkHoldWrRmt_54 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_339) begin
                      cntLkHoldWrRmt_55 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_340) begin
                      cntLkHoldWrRmt_56 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_341) begin
                      cntLkHoldWrRmt_57 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_342) begin
                      cntLkHoldWrRmt_58 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_343) begin
                      cntLkHoldWrRmt_59 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_344) begin
                      cntLkHoldWrRmt_60 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_345) begin
                      cntLkHoldWrRmt_61 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_346) begin
                      cntLkHoldWrRmt_62 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                    if(_zz_347) begin
                      cntLkHoldWrRmt_63 <= _zz_cntLkHoldWrRmt_0_2;
                    end
                  end
                  default : begin
                  end
                endcase
              end
              LockRespType_waiting : begin
                if(_zz_11[0]) begin
                  cntLkWaitRmt_0 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[1]) begin
                  cntLkWaitRmt_1 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[2]) begin
                  cntLkWaitRmt_2 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[3]) begin
                  cntLkWaitRmt_3 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[4]) begin
                  cntLkWaitRmt_4 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[5]) begin
                  cntLkWaitRmt_5 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[6]) begin
                  cntLkWaitRmt_6 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[7]) begin
                  cntLkWaitRmt_7 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[8]) begin
                  cntLkWaitRmt_8 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[9]) begin
                  cntLkWaitRmt_9 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[10]) begin
                  cntLkWaitRmt_10 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[11]) begin
                  cntLkWaitRmt_11 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[12]) begin
                  cntLkWaitRmt_12 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[13]) begin
                  cntLkWaitRmt_13 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[14]) begin
                  cntLkWaitRmt_14 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[15]) begin
                  cntLkWaitRmt_15 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[16]) begin
                  cntLkWaitRmt_16 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[17]) begin
                  cntLkWaitRmt_17 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[18]) begin
                  cntLkWaitRmt_18 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[19]) begin
                  cntLkWaitRmt_19 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[20]) begin
                  cntLkWaitRmt_20 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[21]) begin
                  cntLkWaitRmt_21 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[22]) begin
                  cntLkWaitRmt_22 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[23]) begin
                  cntLkWaitRmt_23 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[24]) begin
                  cntLkWaitRmt_24 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[25]) begin
                  cntLkWaitRmt_25 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[26]) begin
                  cntLkWaitRmt_26 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[27]) begin
                  cntLkWaitRmt_27 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[28]) begin
                  cntLkWaitRmt_28 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[29]) begin
                  cntLkWaitRmt_29 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[30]) begin
                  cntLkWaitRmt_30 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[31]) begin
                  cntLkWaitRmt_31 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[32]) begin
                  cntLkWaitRmt_32 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[33]) begin
                  cntLkWaitRmt_33 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[34]) begin
                  cntLkWaitRmt_34 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[35]) begin
                  cntLkWaitRmt_35 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[36]) begin
                  cntLkWaitRmt_36 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[37]) begin
                  cntLkWaitRmt_37 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[38]) begin
                  cntLkWaitRmt_38 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[39]) begin
                  cntLkWaitRmt_39 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[40]) begin
                  cntLkWaitRmt_40 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[41]) begin
                  cntLkWaitRmt_41 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[42]) begin
                  cntLkWaitRmt_42 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[43]) begin
                  cntLkWaitRmt_43 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[44]) begin
                  cntLkWaitRmt_44 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[45]) begin
                  cntLkWaitRmt_45 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[46]) begin
                  cntLkWaitRmt_46 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[47]) begin
                  cntLkWaitRmt_47 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[48]) begin
                  cntLkWaitRmt_48 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[49]) begin
                  cntLkWaitRmt_49 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[50]) begin
                  cntLkWaitRmt_50 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[51]) begin
                  cntLkWaitRmt_51 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[52]) begin
                  cntLkWaitRmt_52 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[53]) begin
                  cntLkWaitRmt_53 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[54]) begin
                  cntLkWaitRmt_54 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[55]) begin
                  cntLkWaitRmt_55 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[56]) begin
                  cntLkWaitRmt_56 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[57]) begin
                  cntLkWaitRmt_57 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[58]) begin
                  cntLkWaitRmt_58 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[59]) begin
                  cntLkWaitRmt_59 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[60]) begin
                  cntLkWaitRmt_60 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[61]) begin
                  cntLkWaitRmt_61 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[62]) begin
                  cntLkWaitRmt_62 <= _zz_cntLkWaitRmt_0_1;
                end
                if(_zz_11[63]) begin
                  cntLkWaitRmt_63 <= _zz_cntLkWaitRmt_0_1;
                end
              end
              LockRespType_abort : begin
                if(_zz_348[0]) begin
                  rAbort_0 <= 1'b1;
                end
                if(_zz_348[1]) begin
                  rAbort_1 <= 1'b1;
                end
                if(_zz_348[2]) begin
                  rAbort_2 <= 1'b1;
                end
                if(_zz_348[3]) begin
                  rAbort_3 <= 1'b1;
                end
                if(_zz_348[4]) begin
                  rAbort_4 <= 1'b1;
                end
                if(_zz_348[5]) begin
                  rAbort_5 <= 1'b1;
                end
                if(_zz_348[6]) begin
                  rAbort_6 <= 1'b1;
                end
                if(_zz_348[7]) begin
                  rAbort_7 <= 1'b1;
                end
                if(_zz_348[8]) begin
                  rAbort_8 <= 1'b1;
                end
                if(_zz_348[9]) begin
                  rAbort_9 <= 1'b1;
                end
                if(_zz_348[10]) begin
                  rAbort_10 <= 1'b1;
                end
                if(_zz_348[11]) begin
                  rAbort_11 <= 1'b1;
                end
                if(_zz_348[12]) begin
                  rAbort_12 <= 1'b1;
                end
                if(_zz_348[13]) begin
                  rAbort_13 <= 1'b1;
                end
                if(_zz_348[14]) begin
                  rAbort_14 <= 1'b1;
                end
                if(_zz_348[15]) begin
                  rAbort_15 <= 1'b1;
                end
                if(_zz_348[16]) begin
                  rAbort_16 <= 1'b1;
                end
                if(_zz_348[17]) begin
                  rAbort_17 <= 1'b1;
                end
                if(_zz_348[18]) begin
                  rAbort_18 <= 1'b1;
                end
                if(_zz_348[19]) begin
                  rAbort_19 <= 1'b1;
                end
                if(_zz_348[20]) begin
                  rAbort_20 <= 1'b1;
                end
                if(_zz_348[21]) begin
                  rAbort_21 <= 1'b1;
                end
                if(_zz_348[22]) begin
                  rAbort_22 <= 1'b1;
                end
                if(_zz_348[23]) begin
                  rAbort_23 <= 1'b1;
                end
                if(_zz_348[24]) begin
                  rAbort_24 <= 1'b1;
                end
                if(_zz_348[25]) begin
                  rAbort_25 <= 1'b1;
                end
                if(_zz_348[26]) begin
                  rAbort_26 <= 1'b1;
                end
                if(_zz_348[27]) begin
                  rAbort_27 <= 1'b1;
                end
                if(_zz_348[28]) begin
                  rAbort_28 <= 1'b1;
                end
                if(_zz_348[29]) begin
                  rAbort_29 <= 1'b1;
                end
                if(_zz_348[30]) begin
                  rAbort_30 <= 1'b1;
                end
                if(_zz_348[31]) begin
                  rAbort_31 <= 1'b1;
                end
                if(_zz_348[32]) begin
                  rAbort_32 <= 1'b1;
                end
                if(_zz_348[33]) begin
                  rAbort_33 <= 1'b1;
                end
                if(_zz_348[34]) begin
                  rAbort_34 <= 1'b1;
                end
                if(_zz_348[35]) begin
                  rAbort_35 <= 1'b1;
                end
                if(_zz_348[36]) begin
                  rAbort_36 <= 1'b1;
                end
                if(_zz_348[37]) begin
                  rAbort_37 <= 1'b1;
                end
                if(_zz_348[38]) begin
                  rAbort_38 <= 1'b1;
                end
                if(_zz_348[39]) begin
                  rAbort_39 <= 1'b1;
                end
                if(_zz_348[40]) begin
                  rAbort_40 <= 1'b1;
                end
                if(_zz_348[41]) begin
                  rAbort_41 <= 1'b1;
                end
                if(_zz_348[42]) begin
                  rAbort_42 <= 1'b1;
                end
                if(_zz_348[43]) begin
                  rAbort_43 <= 1'b1;
                end
                if(_zz_348[44]) begin
                  rAbort_44 <= 1'b1;
                end
                if(_zz_348[45]) begin
                  rAbort_45 <= 1'b1;
                end
                if(_zz_348[46]) begin
                  rAbort_46 <= 1'b1;
                end
                if(_zz_348[47]) begin
                  rAbort_47 <= 1'b1;
                end
                if(_zz_348[48]) begin
                  rAbort_48 <= 1'b1;
                end
                if(_zz_348[49]) begin
                  rAbort_49 <= 1'b1;
                end
                if(_zz_348[50]) begin
                  rAbort_50 <= 1'b1;
                end
                if(_zz_348[51]) begin
                  rAbort_51 <= 1'b1;
                end
                if(_zz_348[52]) begin
                  rAbort_52 <= 1'b1;
                end
                if(_zz_348[53]) begin
                  rAbort_53 <= 1'b1;
                end
                if(_zz_348[54]) begin
                  rAbort_54 <= 1'b1;
                end
                if(_zz_348[55]) begin
                  rAbort_55 <= 1'b1;
                end
                if(_zz_348[56]) begin
                  rAbort_56 <= 1'b1;
                end
                if(_zz_348[57]) begin
                  rAbort_57 <= 1'b1;
                end
                if(_zz_348[58]) begin
                  rAbort_58 <= 1'b1;
                end
                if(_zz_348[59]) begin
                  rAbort_59 <= 1'b1;
                end
                if(_zz_348[60]) begin
                  rAbort_60 <= 1'b1;
                end
                if(_zz_348[61]) begin
                  rAbort_61 <= 1'b1;
                end
                if(_zz_348[62]) begin
                  rAbort_62 <= 1'b1;
                end
                if(_zz_348[63]) begin
                  rAbort_63 <= 1'b1;
                end
                if(_zz_219) begin
                  cntLkRespRmt_0 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_220) begin
                  cntLkRespRmt_1 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_221) begin
                  cntLkRespRmt_2 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_222) begin
                  cntLkRespRmt_3 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_223) begin
                  cntLkRespRmt_4 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_224) begin
                  cntLkRespRmt_5 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_225) begin
                  cntLkRespRmt_6 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_226) begin
                  cntLkRespRmt_7 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_227) begin
                  cntLkRespRmt_8 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_228) begin
                  cntLkRespRmt_9 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_229) begin
                  cntLkRespRmt_10 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_230) begin
                  cntLkRespRmt_11 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_231) begin
                  cntLkRespRmt_12 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_232) begin
                  cntLkRespRmt_13 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_233) begin
                  cntLkRespRmt_14 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_234) begin
                  cntLkRespRmt_15 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_235) begin
                  cntLkRespRmt_16 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_236) begin
                  cntLkRespRmt_17 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_237) begin
                  cntLkRespRmt_18 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_238) begin
                  cntLkRespRmt_19 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_239) begin
                  cntLkRespRmt_20 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_240) begin
                  cntLkRespRmt_21 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_241) begin
                  cntLkRespRmt_22 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_242) begin
                  cntLkRespRmt_23 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_243) begin
                  cntLkRespRmt_24 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_244) begin
                  cntLkRespRmt_25 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_245) begin
                  cntLkRespRmt_26 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_246) begin
                  cntLkRespRmt_27 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_247) begin
                  cntLkRespRmt_28 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_248) begin
                  cntLkRespRmt_29 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_249) begin
                  cntLkRespRmt_30 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_250) begin
                  cntLkRespRmt_31 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_251) begin
                  cntLkRespRmt_32 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_252) begin
                  cntLkRespRmt_33 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_253) begin
                  cntLkRespRmt_34 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_254) begin
                  cntLkRespRmt_35 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_255) begin
                  cntLkRespRmt_36 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_256) begin
                  cntLkRespRmt_37 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_257) begin
                  cntLkRespRmt_38 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_258) begin
                  cntLkRespRmt_39 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_259) begin
                  cntLkRespRmt_40 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_260) begin
                  cntLkRespRmt_41 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_261) begin
                  cntLkRespRmt_42 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_262) begin
                  cntLkRespRmt_43 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_263) begin
                  cntLkRespRmt_44 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_264) begin
                  cntLkRespRmt_45 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_265) begin
                  cntLkRespRmt_46 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_266) begin
                  cntLkRespRmt_47 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_267) begin
                  cntLkRespRmt_48 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_268) begin
                  cntLkRespRmt_49 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_269) begin
                  cntLkRespRmt_50 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_270) begin
                  cntLkRespRmt_51 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_271) begin
                  cntLkRespRmt_52 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_272) begin
                  cntLkRespRmt_53 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_273) begin
                  cntLkRespRmt_54 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_274) begin
                  cntLkRespRmt_55 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_275) begin
                  cntLkRespRmt_56 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_276) begin
                  cntLkRespRmt_57 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_277) begin
                  cntLkRespRmt_58 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_278) begin
                  cntLkRespRmt_59 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_279) begin
                  cntLkRespRmt_60 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_280) begin
                  cntLkRespRmt_61 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_281) begin
                  cntLkRespRmt_62 <= _zz_cntLkRespRmt_0_2;
                end
                if(_zz_282) begin
                  cntLkRespRmt_63 <= _zz_cntLkRespRmt_0_2;
                end
                io_cntLockDenyRmt <= (io_cntLockDenyRmt + 32'h00000001);
              end
              default : begin
                if(_zz_9[0]) begin
                  cntRlseRespRmt_0 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[1]) begin
                  cntRlseRespRmt_1 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[2]) begin
                  cntRlseRespRmt_2 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[3]) begin
                  cntRlseRespRmt_3 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[4]) begin
                  cntRlseRespRmt_4 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[5]) begin
                  cntRlseRespRmt_5 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[6]) begin
                  cntRlseRespRmt_6 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[7]) begin
                  cntRlseRespRmt_7 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[8]) begin
                  cntRlseRespRmt_8 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[9]) begin
                  cntRlseRespRmt_9 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[10]) begin
                  cntRlseRespRmt_10 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[11]) begin
                  cntRlseRespRmt_11 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[12]) begin
                  cntRlseRespRmt_12 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[13]) begin
                  cntRlseRespRmt_13 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[14]) begin
                  cntRlseRespRmt_14 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[15]) begin
                  cntRlseRespRmt_15 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[16]) begin
                  cntRlseRespRmt_16 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[17]) begin
                  cntRlseRespRmt_17 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[18]) begin
                  cntRlseRespRmt_18 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[19]) begin
                  cntRlseRespRmt_19 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[20]) begin
                  cntRlseRespRmt_20 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[21]) begin
                  cntRlseRespRmt_21 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[22]) begin
                  cntRlseRespRmt_22 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[23]) begin
                  cntRlseRespRmt_23 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[24]) begin
                  cntRlseRespRmt_24 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[25]) begin
                  cntRlseRespRmt_25 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[26]) begin
                  cntRlseRespRmt_26 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[27]) begin
                  cntRlseRespRmt_27 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[28]) begin
                  cntRlseRespRmt_28 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[29]) begin
                  cntRlseRespRmt_29 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[30]) begin
                  cntRlseRespRmt_30 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[31]) begin
                  cntRlseRespRmt_31 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[32]) begin
                  cntRlseRespRmt_32 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[33]) begin
                  cntRlseRespRmt_33 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[34]) begin
                  cntRlseRespRmt_34 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[35]) begin
                  cntRlseRespRmt_35 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[36]) begin
                  cntRlseRespRmt_36 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[37]) begin
                  cntRlseRespRmt_37 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[38]) begin
                  cntRlseRespRmt_38 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[39]) begin
                  cntRlseRespRmt_39 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[40]) begin
                  cntRlseRespRmt_40 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[41]) begin
                  cntRlseRespRmt_41 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[42]) begin
                  cntRlseRespRmt_42 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[43]) begin
                  cntRlseRespRmt_43 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[44]) begin
                  cntRlseRespRmt_44 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[45]) begin
                  cntRlseRespRmt_45 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[46]) begin
                  cntRlseRespRmt_46 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[47]) begin
                  cntRlseRespRmt_47 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[48]) begin
                  cntRlseRespRmt_48 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[49]) begin
                  cntRlseRespRmt_49 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[50]) begin
                  cntRlseRespRmt_50 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[51]) begin
                  cntRlseRespRmt_51 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[52]) begin
                  cntRlseRespRmt_52 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[53]) begin
                  cntRlseRespRmt_53 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[54]) begin
                  cntRlseRespRmt_54 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[55]) begin
                  cntRlseRespRmt_55 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[56]) begin
                  cntRlseRespRmt_56 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[57]) begin
                  cntRlseRespRmt_57 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[58]) begin
                  cntRlseRespRmt_58 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[59]) begin
                  cntRlseRespRmt_59 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[60]) begin
                  cntRlseRespRmt_60 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[61]) begin
                  cntRlseRespRmt_61 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[62]) begin
                  cntRlseRespRmt_62 <= _zz_cntRlseRespRmt_0_1;
                end
                if(_zz_9[63]) begin
                  cntRlseRespRmt_63 <= _zz_cntRlseRespRmt_0_1;
                end
              end
            endcase
          end
        end
        compLkRespRmt_enumDef_RMT_RD_CONSUME : begin
          if(io_rdRmt_fire) begin
            compLkRespRmt_nBeat <= (compLkRespRmt_nBeat + 8'h01);
            if(when_TxnManCS_l315) begin
              compLkRespRmt_nBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
      compTxnCmtLoc_stateReg <= compTxnCmtLoc_stateNext;
      case(compTxnCmtLoc_stateReg)
        compTxnCmtLoc_enumDef_CS_TXN : begin
          if(!when_TxnManCS_l369) begin
            compTxnCmtLoc_curTxnId <= (compTxnCmtLoc_curTxnId + 6'h01);
          end
        end
        compTxnCmtLoc_enumDef_LOCAL_AW : begin
        end
        compTxnCmtLoc_enumDef_LOCAL_W : begin
          if(io_axi_w_fire) begin
            compTxnCmtLoc_nBeat <= (compTxnCmtLoc_nBeat + 8'h01);
            if(io_axi_w_payload_last) begin
              if(_zz_14[0]) begin
                cntCmtReqLoc_0 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[1]) begin
                cntCmtReqLoc_1 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[2]) begin
                cntCmtReqLoc_2 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[3]) begin
                cntCmtReqLoc_3 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[4]) begin
                cntCmtReqLoc_4 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[5]) begin
                cntCmtReqLoc_5 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[6]) begin
                cntCmtReqLoc_6 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[7]) begin
                cntCmtReqLoc_7 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[8]) begin
                cntCmtReqLoc_8 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[9]) begin
                cntCmtReqLoc_9 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[10]) begin
                cntCmtReqLoc_10 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[11]) begin
                cntCmtReqLoc_11 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[12]) begin
                cntCmtReqLoc_12 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[13]) begin
                cntCmtReqLoc_13 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[14]) begin
                cntCmtReqLoc_14 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[15]) begin
                cntCmtReqLoc_15 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[16]) begin
                cntCmtReqLoc_16 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[17]) begin
                cntCmtReqLoc_17 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[18]) begin
                cntCmtReqLoc_18 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[19]) begin
                cntCmtReqLoc_19 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[20]) begin
                cntCmtReqLoc_20 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[21]) begin
                cntCmtReqLoc_21 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[22]) begin
                cntCmtReqLoc_22 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[23]) begin
                cntCmtReqLoc_23 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[24]) begin
                cntCmtReqLoc_24 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[25]) begin
                cntCmtReqLoc_25 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[26]) begin
                cntCmtReqLoc_26 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[27]) begin
                cntCmtReqLoc_27 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[28]) begin
                cntCmtReqLoc_28 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[29]) begin
                cntCmtReqLoc_29 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[30]) begin
                cntCmtReqLoc_30 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[31]) begin
                cntCmtReqLoc_31 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[32]) begin
                cntCmtReqLoc_32 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[33]) begin
                cntCmtReqLoc_33 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[34]) begin
                cntCmtReqLoc_34 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[35]) begin
                cntCmtReqLoc_35 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[36]) begin
                cntCmtReqLoc_36 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[37]) begin
                cntCmtReqLoc_37 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[38]) begin
                cntCmtReqLoc_38 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[39]) begin
                cntCmtReqLoc_39 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[40]) begin
                cntCmtReqLoc_40 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[41]) begin
                cntCmtReqLoc_41 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[42]) begin
                cntCmtReqLoc_42 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[43]) begin
                cntCmtReqLoc_43 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[44]) begin
                cntCmtReqLoc_44 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[45]) begin
                cntCmtReqLoc_45 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[46]) begin
                cntCmtReqLoc_46 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[47]) begin
                cntCmtReqLoc_47 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[48]) begin
                cntCmtReqLoc_48 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[49]) begin
                cntCmtReqLoc_49 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[50]) begin
                cntCmtReqLoc_50 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[51]) begin
                cntCmtReqLoc_51 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[52]) begin
                cntCmtReqLoc_52 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[53]) begin
                cntCmtReqLoc_53 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[54]) begin
                cntCmtReqLoc_54 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[55]) begin
                cntCmtReqLoc_55 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[56]) begin
                cntCmtReqLoc_56 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[57]) begin
                cntCmtReqLoc_57 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[58]) begin
                cntCmtReqLoc_58 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[59]) begin
                cntCmtReqLoc_59 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[60]) begin
                cntCmtReqLoc_60 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[61]) begin
                cntCmtReqLoc_61 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[62]) begin
                cntCmtReqLoc_62 <= _zz_cntCmtReqLoc_0_1;
              end
              if(_zz_14[63]) begin
                cntCmtReqLoc_63 <= _zz_cntCmtReqLoc_0_1;
              end
              compTxnCmtLoc_nBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
      compLkRlseLoc_stateReg <= compLkRlseLoc_stateNext;
      case(compLkRlseLoc_stateReg)
        compLkRlseLoc_enumDef_CS_TXN : begin
          if(!when_TxnManCS_l440) begin
            compLkRlseLoc_curTxnId <= (compLkRlseLoc_curTxnId + 6'h01);
          end
        end
        compLkRlseLoc_enumDef_LK_RLSE : begin
          if(lkReqRlseLoc_fire) begin
            if(_zz_15[0]) begin
              cntRlseReqLoc_0 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[1]) begin
              cntRlseReqLoc_1 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[2]) begin
              cntRlseReqLoc_2 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[3]) begin
              cntRlseReqLoc_3 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[4]) begin
              cntRlseReqLoc_4 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[5]) begin
              cntRlseReqLoc_5 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[6]) begin
              cntRlseReqLoc_6 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[7]) begin
              cntRlseReqLoc_7 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[8]) begin
              cntRlseReqLoc_8 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[9]) begin
              cntRlseReqLoc_9 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[10]) begin
              cntRlseReqLoc_10 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[11]) begin
              cntRlseReqLoc_11 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[12]) begin
              cntRlseReqLoc_12 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[13]) begin
              cntRlseReqLoc_13 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[14]) begin
              cntRlseReqLoc_14 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[15]) begin
              cntRlseReqLoc_15 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[16]) begin
              cntRlseReqLoc_16 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[17]) begin
              cntRlseReqLoc_17 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[18]) begin
              cntRlseReqLoc_18 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[19]) begin
              cntRlseReqLoc_19 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[20]) begin
              cntRlseReqLoc_20 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[21]) begin
              cntRlseReqLoc_21 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[22]) begin
              cntRlseReqLoc_22 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[23]) begin
              cntRlseReqLoc_23 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[24]) begin
              cntRlseReqLoc_24 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[25]) begin
              cntRlseReqLoc_25 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[26]) begin
              cntRlseReqLoc_26 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[27]) begin
              cntRlseReqLoc_27 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[28]) begin
              cntRlseReqLoc_28 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[29]) begin
              cntRlseReqLoc_29 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[30]) begin
              cntRlseReqLoc_30 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[31]) begin
              cntRlseReqLoc_31 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[32]) begin
              cntRlseReqLoc_32 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[33]) begin
              cntRlseReqLoc_33 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[34]) begin
              cntRlseReqLoc_34 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[35]) begin
              cntRlseReqLoc_35 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[36]) begin
              cntRlseReqLoc_36 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[37]) begin
              cntRlseReqLoc_37 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[38]) begin
              cntRlseReqLoc_38 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[39]) begin
              cntRlseReqLoc_39 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[40]) begin
              cntRlseReqLoc_40 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[41]) begin
              cntRlseReqLoc_41 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[42]) begin
              cntRlseReqLoc_42 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[43]) begin
              cntRlseReqLoc_43 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[44]) begin
              cntRlseReqLoc_44 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[45]) begin
              cntRlseReqLoc_45 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[46]) begin
              cntRlseReqLoc_46 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[47]) begin
              cntRlseReqLoc_47 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[48]) begin
              cntRlseReqLoc_48 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[49]) begin
              cntRlseReqLoc_49 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[50]) begin
              cntRlseReqLoc_50 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[51]) begin
              cntRlseReqLoc_51 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[52]) begin
              cntRlseReqLoc_52 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[53]) begin
              cntRlseReqLoc_53 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[54]) begin
              cntRlseReqLoc_54 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[55]) begin
              cntRlseReqLoc_55 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[56]) begin
              cntRlseReqLoc_56 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[57]) begin
              cntRlseReqLoc_57 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[58]) begin
              cntRlseReqLoc_58 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[59]) begin
              cntRlseReqLoc_59 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[60]) begin
              cntRlseReqLoc_60 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[61]) begin
              cntRlseReqLoc_61 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[62]) begin
              cntRlseReqLoc_62 <= _zz_cntRlseReqLoc_0_1;
            end
            if(_zz_15[63]) begin
              cntRlseReqLoc_63 <= _zz_cntRlseReqLoc_0_1;
            end
          end
          if(when_TxnManCS_l456) begin
            if(_zz_349[0]) begin
              cntRlseReqWrLoc_0 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[1]) begin
              cntRlseReqWrLoc_1 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[2]) begin
              cntRlseReqWrLoc_2 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[3]) begin
              cntRlseReqWrLoc_3 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[4]) begin
              cntRlseReqWrLoc_4 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[5]) begin
              cntRlseReqWrLoc_5 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[6]) begin
              cntRlseReqWrLoc_6 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[7]) begin
              cntRlseReqWrLoc_7 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[8]) begin
              cntRlseReqWrLoc_8 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[9]) begin
              cntRlseReqWrLoc_9 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[10]) begin
              cntRlseReqWrLoc_10 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[11]) begin
              cntRlseReqWrLoc_11 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[12]) begin
              cntRlseReqWrLoc_12 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[13]) begin
              cntRlseReqWrLoc_13 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[14]) begin
              cntRlseReqWrLoc_14 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[15]) begin
              cntRlseReqWrLoc_15 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[16]) begin
              cntRlseReqWrLoc_16 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[17]) begin
              cntRlseReqWrLoc_17 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[18]) begin
              cntRlseReqWrLoc_18 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[19]) begin
              cntRlseReqWrLoc_19 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[20]) begin
              cntRlseReqWrLoc_20 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[21]) begin
              cntRlseReqWrLoc_21 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[22]) begin
              cntRlseReqWrLoc_22 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[23]) begin
              cntRlseReqWrLoc_23 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[24]) begin
              cntRlseReqWrLoc_24 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[25]) begin
              cntRlseReqWrLoc_25 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[26]) begin
              cntRlseReqWrLoc_26 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[27]) begin
              cntRlseReqWrLoc_27 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[28]) begin
              cntRlseReqWrLoc_28 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[29]) begin
              cntRlseReqWrLoc_29 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[30]) begin
              cntRlseReqWrLoc_30 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[31]) begin
              cntRlseReqWrLoc_31 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[32]) begin
              cntRlseReqWrLoc_32 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[33]) begin
              cntRlseReqWrLoc_33 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[34]) begin
              cntRlseReqWrLoc_34 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[35]) begin
              cntRlseReqWrLoc_35 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[36]) begin
              cntRlseReqWrLoc_36 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[37]) begin
              cntRlseReqWrLoc_37 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[38]) begin
              cntRlseReqWrLoc_38 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[39]) begin
              cntRlseReqWrLoc_39 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[40]) begin
              cntRlseReqWrLoc_40 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[41]) begin
              cntRlseReqWrLoc_41 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[42]) begin
              cntRlseReqWrLoc_42 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[43]) begin
              cntRlseReqWrLoc_43 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[44]) begin
              cntRlseReqWrLoc_44 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[45]) begin
              cntRlseReqWrLoc_45 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[46]) begin
              cntRlseReqWrLoc_46 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[47]) begin
              cntRlseReqWrLoc_47 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[48]) begin
              cntRlseReqWrLoc_48 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[49]) begin
              cntRlseReqWrLoc_49 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[50]) begin
              cntRlseReqWrLoc_50 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[51]) begin
              cntRlseReqWrLoc_51 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[52]) begin
              cntRlseReqWrLoc_52 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[53]) begin
              cntRlseReqWrLoc_53 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[54]) begin
              cntRlseReqWrLoc_54 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[55]) begin
              cntRlseReqWrLoc_55 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[56]) begin
              cntRlseReqWrLoc_56 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[57]) begin
              cntRlseReqWrLoc_57 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[58]) begin
              cntRlseReqWrLoc_58 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[59]) begin
              cntRlseReqWrLoc_59 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[60]) begin
              cntRlseReqWrLoc_60 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[61]) begin
              cntRlseReqWrLoc_61 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[62]) begin
              cntRlseReqWrLoc_62 <= _zz_cntRlseReqWrLoc_0_1;
            end
            if(_zz_349[63]) begin
              cntRlseReqWrLoc_63 <= _zz_cntRlseReqWrLoc_0_1;
            end
          end
        end
        default : begin
        end
      endcase
      compLkRlseRmt_stateReg <= compLkRlseRmt_stateNext;
      case(compLkRlseRmt_stateReg)
        compLkRlseRmt_enumDef_CS_TXN : begin
          if(!when_TxnManCS_l489) begin
            compLkRlseRmt_curTxnId <= (compLkRlseRmt_curTxnId + 6'h01);
          end
        end
        compLkRlseRmt_enumDef_RMT_LK_RLSE : begin
          if(lkReqRlseRmt_fire) begin
            if(when_TxnManCS_l505) begin
              if(_zz_350[0]) begin
                cntRlseReqWrRmt_0 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[1]) begin
                cntRlseReqWrRmt_1 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[2]) begin
                cntRlseReqWrRmt_2 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[3]) begin
                cntRlseReqWrRmt_3 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[4]) begin
                cntRlseReqWrRmt_4 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[5]) begin
                cntRlseReqWrRmt_5 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[6]) begin
                cntRlseReqWrRmt_6 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[7]) begin
                cntRlseReqWrRmt_7 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[8]) begin
                cntRlseReqWrRmt_8 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[9]) begin
                cntRlseReqWrRmt_9 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[10]) begin
                cntRlseReqWrRmt_10 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[11]) begin
                cntRlseReqWrRmt_11 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[12]) begin
                cntRlseReqWrRmt_12 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[13]) begin
                cntRlseReqWrRmt_13 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[14]) begin
                cntRlseReqWrRmt_14 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[15]) begin
                cntRlseReqWrRmt_15 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[16]) begin
                cntRlseReqWrRmt_16 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[17]) begin
                cntRlseReqWrRmt_17 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[18]) begin
                cntRlseReqWrRmt_18 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[19]) begin
                cntRlseReqWrRmt_19 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[20]) begin
                cntRlseReqWrRmt_20 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[21]) begin
                cntRlseReqWrRmt_21 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[22]) begin
                cntRlseReqWrRmt_22 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[23]) begin
                cntRlseReqWrRmt_23 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[24]) begin
                cntRlseReqWrRmt_24 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[25]) begin
                cntRlseReqWrRmt_25 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[26]) begin
                cntRlseReqWrRmt_26 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[27]) begin
                cntRlseReqWrRmt_27 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[28]) begin
                cntRlseReqWrRmt_28 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[29]) begin
                cntRlseReqWrRmt_29 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[30]) begin
                cntRlseReqWrRmt_30 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[31]) begin
                cntRlseReqWrRmt_31 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[32]) begin
                cntRlseReqWrRmt_32 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[33]) begin
                cntRlseReqWrRmt_33 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[34]) begin
                cntRlseReqWrRmt_34 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[35]) begin
                cntRlseReqWrRmt_35 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[36]) begin
                cntRlseReqWrRmt_36 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[37]) begin
                cntRlseReqWrRmt_37 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[38]) begin
                cntRlseReqWrRmt_38 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[39]) begin
                cntRlseReqWrRmt_39 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[40]) begin
                cntRlseReqWrRmt_40 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[41]) begin
                cntRlseReqWrRmt_41 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[42]) begin
                cntRlseReqWrRmt_42 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[43]) begin
                cntRlseReqWrRmt_43 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[44]) begin
                cntRlseReqWrRmt_44 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[45]) begin
                cntRlseReqWrRmt_45 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[46]) begin
                cntRlseReqWrRmt_46 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[47]) begin
                cntRlseReqWrRmt_47 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[48]) begin
                cntRlseReqWrRmt_48 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[49]) begin
                cntRlseReqWrRmt_49 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[50]) begin
                cntRlseReqWrRmt_50 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[51]) begin
                cntRlseReqWrRmt_51 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[52]) begin
                cntRlseReqWrRmt_52 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[53]) begin
                cntRlseReqWrRmt_53 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[54]) begin
                cntRlseReqWrRmt_54 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[55]) begin
                cntRlseReqWrRmt_55 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[56]) begin
                cntRlseReqWrRmt_56 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[57]) begin
                cntRlseReqWrRmt_57 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[58]) begin
                cntRlseReqWrRmt_58 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[59]) begin
                cntRlseReqWrRmt_59 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[60]) begin
                cntRlseReqWrRmt_60 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[61]) begin
                cntRlseReqWrRmt_61 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[62]) begin
                cntRlseReqWrRmt_62 <= _zz_cntRlseReqWrRmt_0;
              end
              if(_zz_350[63]) begin
                cntRlseReqWrRmt_63 <= _zz_cntRlseReqWrRmt_0;
              end
            end else begin
              if(_zz_17) begin
                cntRlseReqRmt_0 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_18) begin
                cntRlseReqRmt_1 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_19) begin
                cntRlseReqRmt_2 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_20) begin
                cntRlseReqRmt_3 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_21) begin
                cntRlseReqRmt_4 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_22) begin
                cntRlseReqRmt_5 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_23) begin
                cntRlseReqRmt_6 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_24) begin
                cntRlseReqRmt_7 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_25) begin
                cntRlseReqRmt_8 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_26) begin
                cntRlseReqRmt_9 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_27) begin
                cntRlseReqRmt_10 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_28) begin
                cntRlseReqRmt_11 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_29) begin
                cntRlseReqRmt_12 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_30) begin
                cntRlseReqRmt_13 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_31) begin
                cntRlseReqRmt_14 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_32) begin
                cntRlseReqRmt_15 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_33) begin
                cntRlseReqRmt_16 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_34) begin
                cntRlseReqRmt_17 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_35) begin
                cntRlseReqRmt_18 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_36) begin
                cntRlseReqRmt_19 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_37) begin
                cntRlseReqRmt_20 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_38) begin
                cntRlseReqRmt_21 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_39) begin
                cntRlseReqRmt_22 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_40) begin
                cntRlseReqRmt_23 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_41) begin
                cntRlseReqRmt_24 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_42) begin
                cntRlseReqRmt_25 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_43) begin
                cntRlseReqRmt_26 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_44) begin
                cntRlseReqRmt_27 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_45) begin
                cntRlseReqRmt_28 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_46) begin
                cntRlseReqRmt_29 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_47) begin
                cntRlseReqRmt_30 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_48) begin
                cntRlseReqRmt_31 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_49) begin
                cntRlseReqRmt_32 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_50) begin
                cntRlseReqRmt_33 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_51) begin
                cntRlseReqRmt_34 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_52) begin
                cntRlseReqRmt_35 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_53) begin
                cntRlseReqRmt_36 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_54) begin
                cntRlseReqRmt_37 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_55) begin
                cntRlseReqRmt_38 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_56) begin
                cntRlseReqRmt_39 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_57) begin
                cntRlseReqRmt_40 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_58) begin
                cntRlseReqRmt_41 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_59) begin
                cntRlseReqRmt_42 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_60) begin
                cntRlseReqRmt_43 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_61) begin
                cntRlseReqRmt_44 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_62) begin
                cntRlseReqRmt_45 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_63) begin
                cntRlseReqRmt_46 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_64) begin
                cntRlseReqRmt_47 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_65) begin
                cntRlseReqRmt_48 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_66) begin
                cntRlseReqRmt_49 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_67) begin
                cntRlseReqRmt_50 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_68) begin
                cntRlseReqRmt_51 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_69) begin
                cntRlseReqRmt_52 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_70) begin
                cntRlseReqRmt_53 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_71) begin
                cntRlseReqRmt_54 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_72) begin
                cntRlseReqRmt_55 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_73) begin
                cntRlseReqRmt_56 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_74) begin
                cntRlseReqRmt_57 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_75) begin
                cntRlseReqRmt_58 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_76) begin
                cntRlseReqRmt_59 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_77) begin
                cntRlseReqRmt_60 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_78) begin
                cntRlseReqRmt_61 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_79) begin
                cntRlseReqRmt_62 <= _zz_cntRlseReqRmt_0_1;
              end
              if(_zz_80) begin
                cntRlseReqRmt_63 <= _zz_cntRlseReqRmt_0_1;
              end
            end
          end
        end
        compLkRlseRmt_enumDef_RMT_WR : begin
          if(io_wrRmt_fire) begin
            compLkRlseRmt_nBeat <= (compLkRlseRmt_nBeat + 8'h01);
            if(when_TxnManCS_l521) begin
              if(_zz_17) begin
                cntRlseReqRmt_0 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_18) begin
                cntRlseReqRmt_1 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_19) begin
                cntRlseReqRmt_2 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_20) begin
                cntRlseReqRmt_3 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_21) begin
                cntRlseReqRmt_4 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_22) begin
                cntRlseReqRmt_5 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_23) begin
                cntRlseReqRmt_6 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_24) begin
                cntRlseReqRmt_7 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_25) begin
                cntRlseReqRmt_8 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_26) begin
                cntRlseReqRmt_9 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_27) begin
                cntRlseReqRmt_10 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_28) begin
                cntRlseReqRmt_11 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_29) begin
                cntRlseReqRmt_12 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_30) begin
                cntRlseReqRmt_13 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_31) begin
                cntRlseReqRmt_14 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_32) begin
                cntRlseReqRmt_15 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_33) begin
                cntRlseReqRmt_16 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_34) begin
                cntRlseReqRmt_17 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_35) begin
                cntRlseReqRmt_18 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_36) begin
                cntRlseReqRmt_19 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_37) begin
                cntRlseReqRmt_20 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_38) begin
                cntRlseReqRmt_21 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_39) begin
                cntRlseReqRmt_22 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_40) begin
                cntRlseReqRmt_23 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_41) begin
                cntRlseReqRmt_24 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_42) begin
                cntRlseReqRmt_25 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_43) begin
                cntRlseReqRmt_26 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_44) begin
                cntRlseReqRmt_27 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_45) begin
                cntRlseReqRmt_28 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_46) begin
                cntRlseReqRmt_29 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_47) begin
                cntRlseReqRmt_30 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_48) begin
                cntRlseReqRmt_31 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_49) begin
                cntRlseReqRmt_32 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_50) begin
                cntRlseReqRmt_33 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_51) begin
                cntRlseReqRmt_34 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_52) begin
                cntRlseReqRmt_35 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_53) begin
                cntRlseReqRmt_36 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_54) begin
                cntRlseReqRmt_37 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_55) begin
                cntRlseReqRmt_38 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_56) begin
                cntRlseReqRmt_39 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_57) begin
                cntRlseReqRmt_40 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_58) begin
                cntRlseReqRmt_41 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_59) begin
                cntRlseReqRmt_42 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_60) begin
                cntRlseReqRmt_43 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_61) begin
                cntRlseReqRmt_44 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_62) begin
                cntRlseReqRmt_45 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_63) begin
                cntRlseReqRmt_46 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_64) begin
                cntRlseReqRmt_47 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_65) begin
                cntRlseReqRmt_48 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_66) begin
                cntRlseReqRmt_49 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_67) begin
                cntRlseReqRmt_50 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_68) begin
                cntRlseReqRmt_51 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_69) begin
                cntRlseReqRmt_52 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_70) begin
                cntRlseReqRmt_53 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_71) begin
                cntRlseReqRmt_54 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_72) begin
                cntRlseReqRmt_55 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_73) begin
                cntRlseReqRmt_56 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_74) begin
                cntRlseReqRmt_57 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_75) begin
                cntRlseReqRmt_58 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_76) begin
                cntRlseReqRmt_59 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_77) begin
                cntRlseReqRmt_60 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_78) begin
                cntRlseReqRmt_61 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_79) begin
                cntRlseReqRmt_62 <= _zz_cntRlseReqRmt_0_2;
              end
              if(_zz_80) begin
                cntRlseReqRmt_63 <= _zz_cntRlseReqRmt_0_2;
              end
              compLkRlseRmt_nBeat <= 8'h0;
            end
          end
        end
        default : begin
        end
      endcase
      compTimeOut_stateReg <= compTimeOut_stateNext;
      case(compTimeOut_stateReg)
        compTimeOut_enumDef_IDLE : begin
          if(io_start) begin
            cntTimeOut_0 <= 24'h0;
            cntTimeOut_1 <= 24'h0;
            cntTimeOut_2 <= 24'h0;
            cntTimeOut_3 <= 24'h0;
            cntTimeOut_4 <= 24'h0;
            cntTimeOut_5 <= 24'h0;
            cntTimeOut_6 <= 24'h0;
            cntTimeOut_7 <= 24'h0;
            cntTimeOut_8 <= 24'h0;
            cntTimeOut_9 <= 24'h0;
            cntTimeOut_10 <= 24'h0;
            cntTimeOut_11 <= 24'h0;
            cntTimeOut_12 <= 24'h0;
            cntTimeOut_13 <= 24'h0;
            cntTimeOut_14 <= 24'h0;
            cntTimeOut_15 <= 24'h0;
            cntTimeOut_16 <= 24'h0;
            cntTimeOut_17 <= 24'h0;
            cntTimeOut_18 <= 24'h0;
            cntTimeOut_19 <= 24'h0;
            cntTimeOut_20 <= 24'h0;
            cntTimeOut_21 <= 24'h0;
            cntTimeOut_22 <= 24'h0;
            cntTimeOut_23 <= 24'h0;
            cntTimeOut_24 <= 24'h0;
            cntTimeOut_25 <= 24'h0;
            cntTimeOut_26 <= 24'h0;
            cntTimeOut_27 <= 24'h0;
            cntTimeOut_28 <= 24'h0;
            cntTimeOut_29 <= 24'h0;
            cntTimeOut_30 <= 24'h0;
            cntTimeOut_31 <= 24'h0;
            cntTimeOut_32 <= 24'h0;
            cntTimeOut_33 <= 24'h0;
            cntTimeOut_34 <= 24'h0;
            cntTimeOut_35 <= 24'h0;
            cntTimeOut_36 <= 24'h0;
            cntTimeOut_37 <= 24'h0;
            cntTimeOut_38 <= 24'h0;
            cntTimeOut_39 <= 24'h0;
            cntTimeOut_40 <= 24'h0;
            cntTimeOut_41 <= 24'h0;
            cntTimeOut_42 <= 24'h0;
            cntTimeOut_43 <= 24'h0;
            cntTimeOut_44 <= 24'h0;
            cntTimeOut_45 <= 24'h0;
            cntTimeOut_46 <= 24'h0;
            cntTimeOut_47 <= 24'h0;
            cntTimeOut_48 <= 24'h0;
            cntTimeOut_49 <= 24'h0;
            cntTimeOut_50 <= 24'h0;
            cntTimeOut_51 <= 24'h0;
            cntTimeOut_52 <= 24'h0;
            cntTimeOut_53 <= 24'h0;
            cntTimeOut_54 <= 24'h0;
            cntTimeOut_55 <= 24'h0;
            cntTimeOut_56 <= 24'h0;
            cntTimeOut_57 <= 24'h0;
            cntTimeOut_58 <= 24'h0;
            cntTimeOut_59 <= 24'h0;
            cntTimeOut_60 <= 24'h0;
            cntTimeOut_61 <= 24'h0;
            cntTimeOut_62 <= 24'h0;
            cntTimeOut_63 <= 24'h0;
            rTimeOut_0 <= 1'b0;
            rTimeOut_1 <= 1'b0;
            rTimeOut_2 <= 1'b0;
            rTimeOut_3 <= 1'b0;
            rTimeOut_4 <= 1'b0;
            rTimeOut_5 <= 1'b0;
            rTimeOut_6 <= 1'b0;
            rTimeOut_7 <= 1'b0;
            rTimeOut_8 <= 1'b0;
            rTimeOut_9 <= 1'b0;
            rTimeOut_10 <= 1'b0;
            rTimeOut_11 <= 1'b0;
            rTimeOut_12 <= 1'b0;
            rTimeOut_13 <= 1'b0;
            rTimeOut_14 <= 1'b0;
            rTimeOut_15 <= 1'b0;
            rTimeOut_16 <= 1'b0;
            rTimeOut_17 <= 1'b0;
            rTimeOut_18 <= 1'b0;
            rTimeOut_19 <= 1'b0;
            rTimeOut_20 <= 1'b0;
            rTimeOut_21 <= 1'b0;
            rTimeOut_22 <= 1'b0;
            rTimeOut_23 <= 1'b0;
            rTimeOut_24 <= 1'b0;
            rTimeOut_25 <= 1'b0;
            rTimeOut_26 <= 1'b0;
            rTimeOut_27 <= 1'b0;
            rTimeOut_28 <= 1'b0;
            rTimeOut_29 <= 1'b0;
            rTimeOut_30 <= 1'b0;
            rTimeOut_31 <= 1'b0;
            rTimeOut_32 <= 1'b0;
            rTimeOut_33 <= 1'b0;
            rTimeOut_34 <= 1'b0;
            rTimeOut_35 <= 1'b0;
            rTimeOut_36 <= 1'b0;
            rTimeOut_37 <= 1'b0;
            rTimeOut_38 <= 1'b0;
            rTimeOut_39 <= 1'b0;
            rTimeOut_40 <= 1'b0;
            rTimeOut_41 <= 1'b0;
            rTimeOut_42 <= 1'b0;
            rTimeOut_43 <= 1'b0;
            rTimeOut_44 <= 1'b0;
            rTimeOut_45 <= 1'b0;
            rTimeOut_46 <= 1'b0;
            rTimeOut_47 <= 1'b0;
            rTimeOut_48 <= 1'b0;
            rTimeOut_49 <= 1'b0;
            rTimeOut_50 <= 1'b0;
            rTimeOut_51 <= 1'b0;
            rTimeOut_52 <= 1'b0;
            rTimeOut_53 <= 1'b0;
            rTimeOut_54 <= 1'b0;
            rTimeOut_55 <= 1'b0;
            rTimeOut_56 <= 1'b0;
            rTimeOut_57 <= 1'b0;
            rTimeOut_58 <= 1'b0;
            rTimeOut_59 <= 1'b0;
            rTimeOut_60 <= 1'b0;
            rTimeOut_61 <= 1'b0;
            rTimeOut_62 <= 1'b0;
            rTimeOut_63 <= 1'b0;
          end
        end
        compTimeOut_enumDef_COUNT : begin
          if(rReqDone_0) begin
            cntTimeOut_0 <= (cntTimeOut_0 + 24'h000001);
          end
          if(rReqDone_1) begin
            cntTimeOut_1 <= (cntTimeOut_1 + 24'h000001);
          end
          if(rReqDone_2) begin
            cntTimeOut_2 <= (cntTimeOut_2 + 24'h000001);
          end
          if(rReqDone_3) begin
            cntTimeOut_3 <= (cntTimeOut_3 + 24'h000001);
          end
          if(rReqDone_4) begin
            cntTimeOut_4 <= (cntTimeOut_4 + 24'h000001);
          end
          if(rReqDone_5) begin
            cntTimeOut_5 <= (cntTimeOut_5 + 24'h000001);
          end
          if(rReqDone_6) begin
            cntTimeOut_6 <= (cntTimeOut_6 + 24'h000001);
          end
          if(rReqDone_7) begin
            cntTimeOut_7 <= (cntTimeOut_7 + 24'h000001);
          end
          if(rReqDone_8) begin
            cntTimeOut_8 <= (cntTimeOut_8 + 24'h000001);
          end
          if(rReqDone_9) begin
            cntTimeOut_9 <= (cntTimeOut_9 + 24'h000001);
          end
          if(rReqDone_10) begin
            cntTimeOut_10 <= (cntTimeOut_10 + 24'h000001);
          end
          if(rReqDone_11) begin
            cntTimeOut_11 <= (cntTimeOut_11 + 24'h000001);
          end
          if(rReqDone_12) begin
            cntTimeOut_12 <= (cntTimeOut_12 + 24'h000001);
          end
          if(rReqDone_13) begin
            cntTimeOut_13 <= (cntTimeOut_13 + 24'h000001);
          end
          if(rReqDone_14) begin
            cntTimeOut_14 <= (cntTimeOut_14 + 24'h000001);
          end
          if(rReqDone_15) begin
            cntTimeOut_15 <= (cntTimeOut_15 + 24'h000001);
          end
          if(rReqDone_16) begin
            cntTimeOut_16 <= (cntTimeOut_16 + 24'h000001);
          end
          if(rReqDone_17) begin
            cntTimeOut_17 <= (cntTimeOut_17 + 24'h000001);
          end
          if(rReqDone_18) begin
            cntTimeOut_18 <= (cntTimeOut_18 + 24'h000001);
          end
          if(rReqDone_19) begin
            cntTimeOut_19 <= (cntTimeOut_19 + 24'h000001);
          end
          if(rReqDone_20) begin
            cntTimeOut_20 <= (cntTimeOut_20 + 24'h000001);
          end
          if(rReqDone_21) begin
            cntTimeOut_21 <= (cntTimeOut_21 + 24'h000001);
          end
          if(rReqDone_22) begin
            cntTimeOut_22 <= (cntTimeOut_22 + 24'h000001);
          end
          if(rReqDone_23) begin
            cntTimeOut_23 <= (cntTimeOut_23 + 24'h000001);
          end
          if(rReqDone_24) begin
            cntTimeOut_24 <= (cntTimeOut_24 + 24'h000001);
          end
          if(rReqDone_25) begin
            cntTimeOut_25 <= (cntTimeOut_25 + 24'h000001);
          end
          if(rReqDone_26) begin
            cntTimeOut_26 <= (cntTimeOut_26 + 24'h000001);
          end
          if(rReqDone_27) begin
            cntTimeOut_27 <= (cntTimeOut_27 + 24'h000001);
          end
          if(rReqDone_28) begin
            cntTimeOut_28 <= (cntTimeOut_28 + 24'h000001);
          end
          if(rReqDone_29) begin
            cntTimeOut_29 <= (cntTimeOut_29 + 24'h000001);
          end
          if(rReqDone_30) begin
            cntTimeOut_30 <= (cntTimeOut_30 + 24'h000001);
          end
          if(rReqDone_31) begin
            cntTimeOut_31 <= (cntTimeOut_31 + 24'h000001);
          end
          if(rReqDone_32) begin
            cntTimeOut_32 <= (cntTimeOut_32 + 24'h000001);
          end
          if(rReqDone_33) begin
            cntTimeOut_33 <= (cntTimeOut_33 + 24'h000001);
          end
          if(rReqDone_34) begin
            cntTimeOut_34 <= (cntTimeOut_34 + 24'h000001);
          end
          if(rReqDone_35) begin
            cntTimeOut_35 <= (cntTimeOut_35 + 24'h000001);
          end
          if(rReqDone_36) begin
            cntTimeOut_36 <= (cntTimeOut_36 + 24'h000001);
          end
          if(rReqDone_37) begin
            cntTimeOut_37 <= (cntTimeOut_37 + 24'h000001);
          end
          if(rReqDone_38) begin
            cntTimeOut_38 <= (cntTimeOut_38 + 24'h000001);
          end
          if(rReqDone_39) begin
            cntTimeOut_39 <= (cntTimeOut_39 + 24'h000001);
          end
          if(rReqDone_40) begin
            cntTimeOut_40 <= (cntTimeOut_40 + 24'h000001);
          end
          if(rReqDone_41) begin
            cntTimeOut_41 <= (cntTimeOut_41 + 24'h000001);
          end
          if(rReqDone_42) begin
            cntTimeOut_42 <= (cntTimeOut_42 + 24'h000001);
          end
          if(rReqDone_43) begin
            cntTimeOut_43 <= (cntTimeOut_43 + 24'h000001);
          end
          if(rReqDone_44) begin
            cntTimeOut_44 <= (cntTimeOut_44 + 24'h000001);
          end
          if(rReqDone_45) begin
            cntTimeOut_45 <= (cntTimeOut_45 + 24'h000001);
          end
          if(rReqDone_46) begin
            cntTimeOut_46 <= (cntTimeOut_46 + 24'h000001);
          end
          if(rReqDone_47) begin
            cntTimeOut_47 <= (cntTimeOut_47 + 24'h000001);
          end
          if(rReqDone_48) begin
            cntTimeOut_48 <= (cntTimeOut_48 + 24'h000001);
          end
          if(rReqDone_49) begin
            cntTimeOut_49 <= (cntTimeOut_49 + 24'h000001);
          end
          if(rReqDone_50) begin
            cntTimeOut_50 <= (cntTimeOut_50 + 24'h000001);
          end
          if(rReqDone_51) begin
            cntTimeOut_51 <= (cntTimeOut_51 + 24'h000001);
          end
          if(rReqDone_52) begin
            cntTimeOut_52 <= (cntTimeOut_52 + 24'h000001);
          end
          if(rReqDone_53) begin
            cntTimeOut_53 <= (cntTimeOut_53 + 24'h000001);
          end
          if(rReqDone_54) begin
            cntTimeOut_54 <= (cntTimeOut_54 + 24'h000001);
          end
          if(rReqDone_55) begin
            cntTimeOut_55 <= (cntTimeOut_55 + 24'h000001);
          end
          if(rReqDone_56) begin
            cntTimeOut_56 <= (cntTimeOut_56 + 24'h000001);
          end
          if(rReqDone_57) begin
            cntTimeOut_57 <= (cntTimeOut_57 + 24'h000001);
          end
          if(rReqDone_58) begin
            cntTimeOut_58 <= (cntTimeOut_58 + 24'h000001);
          end
          if(rReqDone_59) begin
            cntTimeOut_59 <= (cntTimeOut_59 + 24'h000001);
          end
          if(rReqDone_60) begin
            cntTimeOut_60 <= (cntTimeOut_60 + 24'h000001);
          end
          if(rReqDone_61) begin
            cntTimeOut_61 <= (cntTimeOut_61 + 24'h000001);
          end
          if(rReqDone_62) begin
            cntTimeOut_62 <= (cntTimeOut_62 + 24'h000001);
          end
          if(rReqDone_63) begin
            cntTimeOut_63 <= (cntTimeOut_63 + 24'h000001);
          end
          if(when_TxnManCS_l555) begin
            rTimeOut_0 <= 1'b1;
            rAbort_0 <= 1'b1;
          end
          if(when_TxnManCS_l555_1) begin
            rTimeOut_1 <= 1'b1;
            rAbort_1 <= 1'b1;
          end
          if(when_TxnManCS_l555_2) begin
            rTimeOut_2 <= 1'b1;
            rAbort_2 <= 1'b1;
          end
          if(when_TxnManCS_l555_3) begin
            rTimeOut_3 <= 1'b1;
            rAbort_3 <= 1'b1;
          end
          if(when_TxnManCS_l555_4) begin
            rTimeOut_4 <= 1'b1;
            rAbort_4 <= 1'b1;
          end
          if(when_TxnManCS_l555_5) begin
            rTimeOut_5 <= 1'b1;
            rAbort_5 <= 1'b1;
          end
          if(when_TxnManCS_l555_6) begin
            rTimeOut_6 <= 1'b1;
            rAbort_6 <= 1'b1;
          end
          if(when_TxnManCS_l555_7) begin
            rTimeOut_7 <= 1'b1;
            rAbort_7 <= 1'b1;
          end
          if(when_TxnManCS_l555_8) begin
            rTimeOut_8 <= 1'b1;
            rAbort_8 <= 1'b1;
          end
          if(when_TxnManCS_l555_9) begin
            rTimeOut_9 <= 1'b1;
            rAbort_9 <= 1'b1;
          end
          if(when_TxnManCS_l555_10) begin
            rTimeOut_10 <= 1'b1;
            rAbort_10 <= 1'b1;
          end
          if(when_TxnManCS_l555_11) begin
            rTimeOut_11 <= 1'b1;
            rAbort_11 <= 1'b1;
          end
          if(when_TxnManCS_l555_12) begin
            rTimeOut_12 <= 1'b1;
            rAbort_12 <= 1'b1;
          end
          if(when_TxnManCS_l555_13) begin
            rTimeOut_13 <= 1'b1;
            rAbort_13 <= 1'b1;
          end
          if(when_TxnManCS_l555_14) begin
            rTimeOut_14 <= 1'b1;
            rAbort_14 <= 1'b1;
          end
          if(when_TxnManCS_l555_15) begin
            rTimeOut_15 <= 1'b1;
            rAbort_15 <= 1'b1;
          end
          if(when_TxnManCS_l555_16) begin
            rTimeOut_16 <= 1'b1;
            rAbort_16 <= 1'b1;
          end
          if(when_TxnManCS_l555_17) begin
            rTimeOut_17 <= 1'b1;
            rAbort_17 <= 1'b1;
          end
          if(when_TxnManCS_l555_18) begin
            rTimeOut_18 <= 1'b1;
            rAbort_18 <= 1'b1;
          end
          if(when_TxnManCS_l555_19) begin
            rTimeOut_19 <= 1'b1;
            rAbort_19 <= 1'b1;
          end
          if(when_TxnManCS_l555_20) begin
            rTimeOut_20 <= 1'b1;
            rAbort_20 <= 1'b1;
          end
          if(when_TxnManCS_l555_21) begin
            rTimeOut_21 <= 1'b1;
            rAbort_21 <= 1'b1;
          end
          if(when_TxnManCS_l555_22) begin
            rTimeOut_22 <= 1'b1;
            rAbort_22 <= 1'b1;
          end
          if(when_TxnManCS_l555_23) begin
            rTimeOut_23 <= 1'b1;
            rAbort_23 <= 1'b1;
          end
          if(when_TxnManCS_l555_24) begin
            rTimeOut_24 <= 1'b1;
            rAbort_24 <= 1'b1;
          end
          if(when_TxnManCS_l555_25) begin
            rTimeOut_25 <= 1'b1;
            rAbort_25 <= 1'b1;
          end
          if(when_TxnManCS_l555_26) begin
            rTimeOut_26 <= 1'b1;
            rAbort_26 <= 1'b1;
          end
          if(when_TxnManCS_l555_27) begin
            rTimeOut_27 <= 1'b1;
            rAbort_27 <= 1'b1;
          end
          if(when_TxnManCS_l555_28) begin
            rTimeOut_28 <= 1'b1;
            rAbort_28 <= 1'b1;
          end
          if(when_TxnManCS_l555_29) begin
            rTimeOut_29 <= 1'b1;
            rAbort_29 <= 1'b1;
          end
          if(when_TxnManCS_l555_30) begin
            rTimeOut_30 <= 1'b1;
            rAbort_30 <= 1'b1;
          end
          if(when_TxnManCS_l555_31) begin
            rTimeOut_31 <= 1'b1;
            rAbort_31 <= 1'b1;
          end
          if(when_TxnManCS_l555_32) begin
            rTimeOut_32 <= 1'b1;
            rAbort_32 <= 1'b1;
          end
          if(when_TxnManCS_l555_33) begin
            rTimeOut_33 <= 1'b1;
            rAbort_33 <= 1'b1;
          end
          if(when_TxnManCS_l555_34) begin
            rTimeOut_34 <= 1'b1;
            rAbort_34 <= 1'b1;
          end
          if(when_TxnManCS_l555_35) begin
            rTimeOut_35 <= 1'b1;
            rAbort_35 <= 1'b1;
          end
          if(when_TxnManCS_l555_36) begin
            rTimeOut_36 <= 1'b1;
            rAbort_36 <= 1'b1;
          end
          if(when_TxnManCS_l555_37) begin
            rTimeOut_37 <= 1'b1;
            rAbort_37 <= 1'b1;
          end
          if(when_TxnManCS_l555_38) begin
            rTimeOut_38 <= 1'b1;
            rAbort_38 <= 1'b1;
          end
          if(when_TxnManCS_l555_39) begin
            rTimeOut_39 <= 1'b1;
            rAbort_39 <= 1'b1;
          end
          if(when_TxnManCS_l555_40) begin
            rTimeOut_40 <= 1'b1;
            rAbort_40 <= 1'b1;
          end
          if(when_TxnManCS_l555_41) begin
            rTimeOut_41 <= 1'b1;
            rAbort_41 <= 1'b1;
          end
          if(when_TxnManCS_l555_42) begin
            rTimeOut_42 <= 1'b1;
            rAbort_42 <= 1'b1;
          end
          if(when_TxnManCS_l555_43) begin
            rTimeOut_43 <= 1'b1;
            rAbort_43 <= 1'b1;
          end
          if(when_TxnManCS_l555_44) begin
            rTimeOut_44 <= 1'b1;
            rAbort_44 <= 1'b1;
          end
          if(when_TxnManCS_l555_45) begin
            rTimeOut_45 <= 1'b1;
            rAbort_45 <= 1'b1;
          end
          if(when_TxnManCS_l555_46) begin
            rTimeOut_46 <= 1'b1;
            rAbort_46 <= 1'b1;
          end
          if(when_TxnManCS_l555_47) begin
            rTimeOut_47 <= 1'b1;
            rAbort_47 <= 1'b1;
          end
          if(when_TxnManCS_l555_48) begin
            rTimeOut_48 <= 1'b1;
            rAbort_48 <= 1'b1;
          end
          if(when_TxnManCS_l555_49) begin
            rTimeOut_49 <= 1'b1;
            rAbort_49 <= 1'b1;
          end
          if(when_TxnManCS_l555_50) begin
            rTimeOut_50 <= 1'b1;
            rAbort_50 <= 1'b1;
          end
          if(when_TxnManCS_l555_51) begin
            rTimeOut_51 <= 1'b1;
            rAbort_51 <= 1'b1;
          end
          if(when_TxnManCS_l555_52) begin
            rTimeOut_52 <= 1'b1;
            rAbort_52 <= 1'b1;
          end
          if(when_TxnManCS_l555_53) begin
            rTimeOut_53 <= 1'b1;
            rAbort_53 <= 1'b1;
          end
          if(when_TxnManCS_l555_54) begin
            rTimeOut_54 <= 1'b1;
            rAbort_54 <= 1'b1;
          end
          if(when_TxnManCS_l555_55) begin
            rTimeOut_55 <= 1'b1;
            rAbort_55 <= 1'b1;
          end
          if(when_TxnManCS_l555_56) begin
            rTimeOut_56 <= 1'b1;
            rAbort_56 <= 1'b1;
          end
          if(when_TxnManCS_l555_57) begin
            rTimeOut_57 <= 1'b1;
            rAbort_57 <= 1'b1;
          end
          if(when_TxnManCS_l555_58) begin
            rTimeOut_58 <= 1'b1;
            rAbort_58 <= 1'b1;
          end
          if(when_TxnManCS_l555_59) begin
            rTimeOut_59 <= 1'b1;
            rAbort_59 <= 1'b1;
          end
          if(when_TxnManCS_l555_60) begin
            rTimeOut_60 <= 1'b1;
            rAbort_60 <= 1'b1;
          end
          if(when_TxnManCS_l555_61) begin
            rTimeOut_61 <= 1'b1;
            rAbort_61 <= 1'b1;
          end
          if(when_TxnManCS_l555_62) begin
            rTimeOut_62 <= 1'b1;
            rAbort_62 <= 1'b1;
          end
          if(when_TxnManCS_l555_63) begin
            rTimeOut_63 <= 1'b1;
            rAbort_63 <= 1'b1;
          end
        end
        default : begin
        end
      endcase
      compLoadTxn_stateReg <= compLoadTxn_stateNext;
      case(compLoadTxn_stateReg)
        compLoadTxn_enumDef_IDLE : begin
          if(io_start) begin
            compLoadTxn_curTxnId <= 6'h0;
            compLoadTxn_cntTxn <= 32'h0;
          end
        end
        compLoadTxn_enumDef_CS_TXN : begin
          if(!when_TxnManCS_l621) begin
            compLoadTxn_curTxnId <= (compLoadTxn_curTxnId + 6'h01);
          end
        end
        compLoadTxn_enumDef_RD_CMDAXI : begin
          if(io_cmdAxi_ar_fire) begin
            compLoadTxn_rTxnMemLd <= 1'b0;
          end
        end
        compLoadTxn_enumDef_LD_TXN : begin
          if(io_cmdAxi_r_fire_2) begin
            compLoadTxn_rTxnMemLd <= 1'b1;
          end
          if(compLoadTxn_cntTxnWordInLine_willOverflow) begin
            compLoadTxn_rTxnMemLd <= 1'b0;
          end
          if(compLoadTxn_cntTxnWord_willOverflow) begin
            if(_zz_354[0]) begin
              cntLkReqLoc_0 <= 6'h0;
            end
            if(_zz_354[1]) begin
              cntLkReqLoc_1 <= 6'h0;
            end
            if(_zz_354[2]) begin
              cntLkReqLoc_2 <= 6'h0;
            end
            if(_zz_354[3]) begin
              cntLkReqLoc_3 <= 6'h0;
            end
            if(_zz_354[4]) begin
              cntLkReqLoc_4 <= 6'h0;
            end
            if(_zz_354[5]) begin
              cntLkReqLoc_5 <= 6'h0;
            end
            if(_zz_354[6]) begin
              cntLkReqLoc_6 <= 6'h0;
            end
            if(_zz_354[7]) begin
              cntLkReqLoc_7 <= 6'h0;
            end
            if(_zz_354[8]) begin
              cntLkReqLoc_8 <= 6'h0;
            end
            if(_zz_354[9]) begin
              cntLkReqLoc_9 <= 6'h0;
            end
            if(_zz_354[10]) begin
              cntLkReqLoc_10 <= 6'h0;
            end
            if(_zz_354[11]) begin
              cntLkReqLoc_11 <= 6'h0;
            end
            if(_zz_354[12]) begin
              cntLkReqLoc_12 <= 6'h0;
            end
            if(_zz_354[13]) begin
              cntLkReqLoc_13 <= 6'h0;
            end
            if(_zz_354[14]) begin
              cntLkReqLoc_14 <= 6'h0;
            end
            if(_zz_354[15]) begin
              cntLkReqLoc_15 <= 6'h0;
            end
            if(_zz_354[16]) begin
              cntLkReqLoc_16 <= 6'h0;
            end
            if(_zz_354[17]) begin
              cntLkReqLoc_17 <= 6'h0;
            end
            if(_zz_354[18]) begin
              cntLkReqLoc_18 <= 6'h0;
            end
            if(_zz_354[19]) begin
              cntLkReqLoc_19 <= 6'h0;
            end
            if(_zz_354[20]) begin
              cntLkReqLoc_20 <= 6'h0;
            end
            if(_zz_354[21]) begin
              cntLkReqLoc_21 <= 6'h0;
            end
            if(_zz_354[22]) begin
              cntLkReqLoc_22 <= 6'h0;
            end
            if(_zz_354[23]) begin
              cntLkReqLoc_23 <= 6'h0;
            end
            if(_zz_354[24]) begin
              cntLkReqLoc_24 <= 6'h0;
            end
            if(_zz_354[25]) begin
              cntLkReqLoc_25 <= 6'h0;
            end
            if(_zz_354[26]) begin
              cntLkReqLoc_26 <= 6'h0;
            end
            if(_zz_354[27]) begin
              cntLkReqLoc_27 <= 6'h0;
            end
            if(_zz_354[28]) begin
              cntLkReqLoc_28 <= 6'h0;
            end
            if(_zz_354[29]) begin
              cntLkReqLoc_29 <= 6'h0;
            end
            if(_zz_354[30]) begin
              cntLkReqLoc_30 <= 6'h0;
            end
            if(_zz_354[31]) begin
              cntLkReqLoc_31 <= 6'h0;
            end
            if(_zz_354[32]) begin
              cntLkReqLoc_32 <= 6'h0;
            end
            if(_zz_354[33]) begin
              cntLkReqLoc_33 <= 6'h0;
            end
            if(_zz_354[34]) begin
              cntLkReqLoc_34 <= 6'h0;
            end
            if(_zz_354[35]) begin
              cntLkReqLoc_35 <= 6'h0;
            end
            if(_zz_354[36]) begin
              cntLkReqLoc_36 <= 6'h0;
            end
            if(_zz_354[37]) begin
              cntLkReqLoc_37 <= 6'h0;
            end
            if(_zz_354[38]) begin
              cntLkReqLoc_38 <= 6'h0;
            end
            if(_zz_354[39]) begin
              cntLkReqLoc_39 <= 6'h0;
            end
            if(_zz_354[40]) begin
              cntLkReqLoc_40 <= 6'h0;
            end
            if(_zz_354[41]) begin
              cntLkReqLoc_41 <= 6'h0;
            end
            if(_zz_354[42]) begin
              cntLkReqLoc_42 <= 6'h0;
            end
            if(_zz_354[43]) begin
              cntLkReqLoc_43 <= 6'h0;
            end
            if(_zz_354[44]) begin
              cntLkReqLoc_44 <= 6'h0;
            end
            if(_zz_354[45]) begin
              cntLkReqLoc_45 <= 6'h0;
            end
            if(_zz_354[46]) begin
              cntLkReqLoc_46 <= 6'h0;
            end
            if(_zz_354[47]) begin
              cntLkReqLoc_47 <= 6'h0;
            end
            if(_zz_354[48]) begin
              cntLkReqLoc_48 <= 6'h0;
            end
            if(_zz_354[49]) begin
              cntLkReqLoc_49 <= 6'h0;
            end
            if(_zz_354[50]) begin
              cntLkReqLoc_50 <= 6'h0;
            end
            if(_zz_354[51]) begin
              cntLkReqLoc_51 <= 6'h0;
            end
            if(_zz_354[52]) begin
              cntLkReqLoc_52 <= 6'h0;
            end
            if(_zz_354[53]) begin
              cntLkReqLoc_53 <= 6'h0;
            end
            if(_zz_354[54]) begin
              cntLkReqLoc_54 <= 6'h0;
            end
            if(_zz_354[55]) begin
              cntLkReqLoc_55 <= 6'h0;
            end
            if(_zz_354[56]) begin
              cntLkReqLoc_56 <= 6'h0;
            end
            if(_zz_354[57]) begin
              cntLkReqLoc_57 <= 6'h0;
            end
            if(_zz_354[58]) begin
              cntLkReqLoc_58 <= 6'h0;
            end
            if(_zz_354[59]) begin
              cntLkReqLoc_59 <= 6'h0;
            end
            if(_zz_354[60]) begin
              cntLkReqLoc_60 <= 6'h0;
            end
            if(_zz_354[61]) begin
              cntLkReqLoc_61 <= 6'h0;
            end
            if(_zz_354[62]) begin
              cntLkReqLoc_62 <= 6'h0;
            end
            if(_zz_354[63]) begin
              cntLkReqLoc_63 <= 6'h0;
            end
            if(_zz_355[0]) begin
              cntLkReqRmt_0 <= 6'h0;
            end
            if(_zz_355[1]) begin
              cntLkReqRmt_1 <= 6'h0;
            end
            if(_zz_355[2]) begin
              cntLkReqRmt_2 <= 6'h0;
            end
            if(_zz_355[3]) begin
              cntLkReqRmt_3 <= 6'h0;
            end
            if(_zz_355[4]) begin
              cntLkReqRmt_4 <= 6'h0;
            end
            if(_zz_355[5]) begin
              cntLkReqRmt_5 <= 6'h0;
            end
            if(_zz_355[6]) begin
              cntLkReqRmt_6 <= 6'h0;
            end
            if(_zz_355[7]) begin
              cntLkReqRmt_7 <= 6'h0;
            end
            if(_zz_355[8]) begin
              cntLkReqRmt_8 <= 6'h0;
            end
            if(_zz_355[9]) begin
              cntLkReqRmt_9 <= 6'h0;
            end
            if(_zz_355[10]) begin
              cntLkReqRmt_10 <= 6'h0;
            end
            if(_zz_355[11]) begin
              cntLkReqRmt_11 <= 6'h0;
            end
            if(_zz_355[12]) begin
              cntLkReqRmt_12 <= 6'h0;
            end
            if(_zz_355[13]) begin
              cntLkReqRmt_13 <= 6'h0;
            end
            if(_zz_355[14]) begin
              cntLkReqRmt_14 <= 6'h0;
            end
            if(_zz_355[15]) begin
              cntLkReqRmt_15 <= 6'h0;
            end
            if(_zz_355[16]) begin
              cntLkReqRmt_16 <= 6'h0;
            end
            if(_zz_355[17]) begin
              cntLkReqRmt_17 <= 6'h0;
            end
            if(_zz_355[18]) begin
              cntLkReqRmt_18 <= 6'h0;
            end
            if(_zz_355[19]) begin
              cntLkReqRmt_19 <= 6'h0;
            end
            if(_zz_355[20]) begin
              cntLkReqRmt_20 <= 6'h0;
            end
            if(_zz_355[21]) begin
              cntLkReqRmt_21 <= 6'h0;
            end
            if(_zz_355[22]) begin
              cntLkReqRmt_22 <= 6'h0;
            end
            if(_zz_355[23]) begin
              cntLkReqRmt_23 <= 6'h0;
            end
            if(_zz_355[24]) begin
              cntLkReqRmt_24 <= 6'h0;
            end
            if(_zz_355[25]) begin
              cntLkReqRmt_25 <= 6'h0;
            end
            if(_zz_355[26]) begin
              cntLkReqRmt_26 <= 6'h0;
            end
            if(_zz_355[27]) begin
              cntLkReqRmt_27 <= 6'h0;
            end
            if(_zz_355[28]) begin
              cntLkReqRmt_28 <= 6'h0;
            end
            if(_zz_355[29]) begin
              cntLkReqRmt_29 <= 6'h0;
            end
            if(_zz_355[30]) begin
              cntLkReqRmt_30 <= 6'h0;
            end
            if(_zz_355[31]) begin
              cntLkReqRmt_31 <= 6'h0;
            end
            if(_zz_355[32]) begin
              cntLkReqRmt_32 <= 6'h0;
            end
            if(_zz_355[33]) begin
              cntLkReqRmt_33 <= 6'h0;
            end
            if(_zz_355[34]) begin
              cntLkReqRmt_34 <= 6'h0;
            end
            if(_zz_355[35]) begin
              cntLkReqRmt_35 <= 6'h0;
            end
            if(_zz_355[36]) begin
              cntLkReqRmt_36 <= 6'h0;
            end
            if(_zz_355[37]) begin
              cntLkReqRmt_37 <= 6'h0;
            end
            if(_zz_355[38]) begin
              cntLkReqRmt_38 <= 6'h0;
            end
            if(_zz_355[39]) begin
              cntLkReqRmt_39 <= 6'h0;
            end
            if(_zz_355[40]) begin
              cntLkReqRmt_40 <= 6'h0;
            end
            if(_zz_355[41]) begin
              cntLkReqRmt_41 <= 6'h0;
            end
            if(_zz_355[42]) begin
              cntLkReqRmt_42 <= 6'h0;
            end
            if(_zz_355[43]) begin
              cntLkReqRmt_43 <= 6'h0;
            end
            if(_zz_355[44]) begin
              cntLkReqRmt_44 <= 6'h0;
            end
            if(_zz_355[45]) begin
              cntLkReqRmt_45 <= 6'h0;
            end
            if(_zz_355[46]) begin
              cntLkReqRmt_46 <= 6'h0;
            end
            if(_zz_355[47]) begin
              cntLkReqRmt_47 <= 6'h0;
            end
            if(_zz_355[48]) begin
              cntLkReqRmt_48 <= 6'h0;
            end
            if(_zz_355[49]) begin
              cntLkReqRmt_49 <= 6'h0;
            end
            if(_zz_355[50]) begin
              cntLkReqRmt_50 <= 6'h0;
            end
            if(_zz_355[51]) begin
              cntLkReqRmt_51 <= 6'h0;
            end
            if(_zz_355[52]) begin
              cntLkReqRmt_52 <= 6'h0;
            end
            if(_zz_355[53]) begin
              cntLkReqRmt_53 <= 6'h0;
            end
            if(_zz_355[54]) begin
              cntLkReqRmt_54 <= 6'h0;
            end
            if(_zz_355[55]) begin
              cntLkReqRmt_55 <= 6'h0;
            end
            if(_zz_355[56]) begin
              cntLkReqRmt_56 <= 6'h0;
            end
            if(_zz_355[57]) begin
              cntLkReqRmt_57 <= 6'h0;
            end
            if(_zz_355[58]) begin
              cntLkReqRmt_58 <= 6'h0;
            end
            if(_zz_355[59]) begin
              cntLkReqRmt_59 <= 6'h0;
            end
            if(_zz_355[60]) begin
              cntLkReqRmt_60 <= 6'h0;
            end
            if(_zz_355[61]) begin
              cntLkReqRmt_61 <= 6'h0;
            end
            if(_zz_355[62]) begin
              cntLkReqRmt_62 <= 6'h0;
            end
            if(_zz_355[63]) begin
              cntLkReqRmt_63 <= 6'h0;
            end
            if(_zz_356[0]) begin
              cntLkRespLoc_0 <= 6'h0;
            end
            if(_zz_356[1]) begin
              cntLkRespLoc_1 <= 6'h0;
            end
            if(_zz_356[2]) begin
              cntLkRespLoc_2 <= 6'h0;
            end
            if(_zz_356[3]) begin
              cntLkRespLoc_3 <= 6'h0;
            end
            if(_zz_356[4]) begin
              cntLkRespLoc_4 <= 6'h0;
            end
            if(_zz_356[5]) begin
              cntLkRespLoc_5 <= 6'h0;
            end
            if(_zz_356[6]) begin
              cntLkRespLoc_6 <= 6'h0;
            end
            if(_zz_356[7]) begin
              cntLkRespLoc_7 <= 6'h0;
            end
            if(_zz_356[8]) begin
              cntLkRespLoc_8 <= 6'h0;
            end
            if(_zz_356[9]) begin
              cntLkRespLoc_9 <= 6'h0;
            end
            if(_zz_356[10]) begin
              cntLkRespLoc_10 <= 6'h0;
            end
            if(_zz_356[11]) begin
              cntLkRespLoc_11 <= 6'h0;
            end
            if(_zz_356[12]) begin
              cntLkRespLoc_12 <= 6'h0;
            end
            if(_zz_356[13]) begin
              cntLkRespLoc_13 <= 6'h0;
            end
            if(_zz_356[14]) begin
              cntLkRespLoc_14 <= 6'h0;
            end
            if(_zz_356[15]) begin
              cntLkRespLoc_15 <= 6'h0;
            end
            if(_zz_356[16]) begin
              cntLkRespLoc_16 <= 6'h0;
            end
            if(_zz_356[17]) begin
              cntLkRespLoc_17 <= 6'h0;
            end
            if(_zz_356[18]) begin
              cntLkRespLoc_18 <= 6'h0;
            end
            if(_zz_356[19]) begin
              cntLkRespLoc_19 <= 6'h0;
            end
            if(_zz_356[20]) begin
              cntLkRespLoc_20 <= 6'h0;
            end
            if(_zz_356[21]) begin
              cntLkRespLoc_21 <= 6'h0;
            end
            if(_zz_356[22]) begin
              cntLkRespLoc_22 <= 6'h0;
            end
            if(_zz_356[23]) begin
              cntLkRespLoc_23 <= 6'h0;
            end
            if(_zz_356[24]) begin
              cntLkRespLoc_24 <= 6'h0;
            end
            if(_zz_356[25]) begin
              cntLkRespLoc_25 <= 6'h0;
            end
            if(_zz_356[26]) begin
              cntLkRespLoc_26 <= 6'h0;
            end
            if(_zz_356[27]) begin
              cntLkRespLoc_27 <= 6'h0;
            end
            if(_zz_356[28]) begin
              cntLkRespLoc_28 <= 6'h0;
            end
            if(_zz_356[29]) begin
              cntLkRespLoc_29 <= 6'h0;
            end
            if(_zz_356[30]) begin
              cntLkRespLoc_30 <= 6'h0;
            end
            if(_zz_356[31]) begin
              cntLkRespLoc_31 <= 6'h0;
            end
            if(_zz_356[32]) begin
              cntLkRespLoc_32 <= 6'h0;
            end
            if(_zz_356[33]) begin
              cntLkRespLoc_33 <= 6'h0;
            end
            if(_zz_356[34]) begin
              cntLkRespLoc_34 <= 6'h0;
            end
            if(_zz_356[35]) begin
              cntLkRespLoc_35 <= 6'h0;
            end
            if(_zz_356[36]) begin
              cntLkRespLoc_36 <= 6'h0;
            end
            if(_zz_356[37]) begin
              cntLkRespLoc_37 <= 6'h0;
            end
            if(_zz_356[38]) begin
              cntLkRespLoc_38 <= 6'h0;
            end
            if(_zz_356[39]) begin
              cntLkRespLoc_39 <= 6'h0;
            end
            if(_zz_356[40]) begin
              cntLkRespLoc_40 <= 6'h0;
            end
            if(_zz_356[41]) begin
              cntLkRespLoc_41 <= 6'h0;
            end
            if(_zz_356[42]) begin
              cntLkRespLoc_42 <= 6'h0;
            end
            if(_zz_356[43]) begin
              cntLkRespLoc_43 <= 6'h0;
            end
            if(_zz_356[44]) begin
              cntLkRespLoc_44 <= 6'h0;
            end
            if(_zz_356[45]) begin
              cntLkRespLoc_45 <= 6'h0;
            end
            if(_zz_356[46]) begin
              cntLkRespLoc_46 <= 6'h0;
            end
            if(_zz_356[47]) begin
              cntLkRespLoc_47 <= 6'h0;
            end
            if(_zz_356[48]) begin
              cntLkRespLoc_48 <= 6'h0;
            end
            if(_zz_356[49]) begin
              cntLkRespLoc_49 <= 6'h0;
            end
            if(_zz_356[50]) begin
              cntLkRespLoc_50 <= 6'h0;
            end
            if(_zz_356[51]) begin
              cntLkRespLoc_51 <= 6'h0;
            end
            if(_zz_356[52]) begin
              cntLkRespLoc_52 <= 6'h0;
            end
            if(_zz_356[53]) begin
              cntLkRespLoc_53 <= 6'h0;
            end
            if(_zz_356[54]) begin
              cntLkRespLoc_54 <= 6'h0;
            end
            if(_zz_356[55]) begin
              cntLkRespLoc_55 <= 6'h0;
            end
            if(_zz_356[56]) begin
              cntLkRespLoc_56 <= 6'h0;
            end
            if(_zz_356[57]) begin
              cntLkRespLoc_57 <= 6'h0;
            end
            if(_zz_356[58]) begin
              cntLkRespLoc_58 <= 6'h0;
            end
            if(_zz_356[59]) begin
              cntLkRespLoc_59 <= 6'h0;
            end
            if(_zz_356[60]) begin
              cntLkRespLoc_60 <= 6'h0;
            end
            if(_zz_356[61]) begin
              cntLkRespLoc_61 <= 6'h0;
            end
            if(_zz_356[62]) begin
              cntLkRespLoc_62 <= 6'h0;
            end
            if(_zz_356[63]) begin
              cntLkRespLoc_63 <= 6'h0;
            end
            if(_zz_357[0]) begin
              cntLkRespRmt_0 <= 6'h0;
            end
            if(_zz_357[1]) begin
              cntLkRespRmt_1 <= 6'h0;
            end
            if(_zz_357[2]) begin
              cntLkRespRmt_2 <= 6'h0;
            end
            if(_zz_357[3]) begin
              cntLkRespRmt_3 <= 6'h0;
            end
            if(_zz_357[4]) begin
              cntLkRespRmt_4 <= 6'h0;
            end
            if(_zz_357[5]) begin
              cntLkRespRmt_5 <= 6'h0;
            end
            if(_zz_357[6]) begin
              cntLkRespRmt_6 <= 6'h0;
            end
            if(_zz_357[7]) begin
              cntLkRespRmt_7 <= 6'h0;
            end
            if(_zz_357[8]) begin
              cntLkRespRmt_8 <= 6'h0;
            end
            if(_zz_357[9]) begin
              cntLkRespRmt_9 <= 6'h0;
            end
            if(_zz_357[10]) begin
              cntLkRespRmt_10 <= 6'h0;
            end
            if(_zz_357[11]) begin
              cntLkRespRmt_11 <= 6'h0;
            end
            if(_zz_357[12]) begin
              cntLkRespRmt_12 <= 6'h0;
            end
            if(_zz_357[13]) begin
              cntLkRespRmt_13 <= 6'h0;
            end
            if(_zz_357[14]) begin
              cntLkRespRmt_14 <= 6'h0;
            end
            if(_zz_357[15]) begin
              cntLkRespRmt_15 <= 6'h0;
            end
            if(_zz_357[16]) begin
              cntLkRespRmt_16 <= 6'h0;
            end
            if(_zz_357[17]) begin
              cntLkRespRmt_17 <= 6'h0;
            end
            if(_zz_357[18]) begin
              cntLkRespRmt_18 <= 6'h0;
            end
            if(_zz_357[19]) begin
              cntLkRespRmt_19 <= 6'h0;
            end
            if(_zz_357[20]) begin
              cntLkRespRmt_20 <= 6'h0;
            end
            if(_zz_357[21]) begin
              cntLkRespRmt_21 <= 6'h0;
            end
            if(_zz_357[22]) begin
              cntLkRespRmt_22 <= 6'h0;
            end
            if(_zz_357[23]) begin
              cntLkRespRmt_23 <= 6'h0;
            end
            if(_zz_357[24]) begin
              cntLkRespRmt_24 <= 6'h0;
            end
            if(_zz_357[25]) begin
              cntLkRespRmt_25 <= 6'h0;
            end
            if(_zz_357[26]) begin
              cntLkRespRmt_26 <= 6'h0;
            end
            if(_zz_357[27]) begin
              cntLkRespRmt_27 <= 6'h0;
            end
            if(_zz_357[28]) begin
              cntLkRespRmt_28 <= 6'h0;
            end
            if(_zz_357[29]) begin
              cntLkRespRmt_29 <= 6'h0;
            end
            if(_zz_357[30]) begin
              cntLkRespRmt_30 <= 6'h0;
            end
            if(_zz_357[31]) begin
              cntLkRespRmt_31 <= 6'h0;
            end
            if(_zz_357[32]) begin
              cntLkRespRmt_32 <= 6'h0;
            end
            if(_zz_357[33]) begin
              cntLkRespRmt_33 <= 6'h0;
            end
            if(_zz_357[34]) begin
              cntLkRespRmt_34 <= 6'h0;
            end
            if(_zz_357[35]) begin
              cntLkRespRmt_35 <= 6'h0;
            end
            if(_zz_357[36]) begin
              cntLkRespRmt_36 <= 6'h0;
            end
            if(_zz_357[37]) begin
              cntLkRespRmt_37 <= 6'h0;
            end
            if(_zz_357[38]) begin
              cntLkRespRmt_38 <= 6'h0;
            end
            if(_zz_357[39]) begin
              cntLkRespRmt_39 <= 6'h0;
            end
            if(_zz_357[40]) begin
              cntLkRespRmt_40 <= 6'h0;
            end
            if(_zz_357[41]) begin
              cntLkRespRmt_41 <= 6'h0;
            end
            if(_zz_357[42]) begin
              cntLkRespRmt_42 <= 6'h0;
            end
            if(_zz_357[43]) begin
              cntLkRespRmt_43 <= 6'h0;
            end
            if(_zz_357[44]) begin
              cntLkRespRmt_44 <= 6'h0;
            end
            if(_zz_357[45]) begin
              cntLkRespRmt_45 <= 6'h0;
            end
            if(_zz_357[46]) begin
              cntLkRespRmt_46 <= 6'h0;
            end
            if(_zz_357[47]) begin
              cntLkRespRmt_47 <= 6'h0;
            end
            if(_zz_357[48]) begin
              cntLkRespRmt_48 <= 6'h0;
            end
            if(_zz_357[49]) begin
              cntLkRespRmt_49 <= 6'h0;
            end
            if(_zz_357[50]) begin
              cntLkRespRmt_50 <= 6'h0;
            end
            if(_zz_357[51]) begin
              cntLkRespRmt_51 <= 6'h0;
            end
            if(_zz_357[52]) begin
              cntLkRespRmt_52 <= 6'h0;
            end
            if(_zz_357[53]) begin
              cntLkRespRmt_53 <= 6'h0;
            end
            if(_zz_357[54]) begin
              cntLkRespRmt_54 <= 6'h0;
            end
            if(_zz_357[55]) begin
              cntLkRespRmt_55 <= 6'h0;
            end
            if(_zz_357[56]) begin
              cntLkRespRmt_56 <= 6'h0;
            end
            if(_zz_357[57]) begin
              cntLkRespRmt_57 <= 6'h0;
            end
            if(_zz_357[58]) begin
              cntLkRespRmt_58 <= 6'h0;
            end
            if(_zz_357[59]) begin
              cntLkRespRmt_59 <= 6'h0;
            end
            if(_zz_357[60]) begin
              cntLkRespRmt_60 <= 6'h0;
            end
            if(_zz_357[61]) begin
              cntLkRespRmt_61 <= 6'h0;
            end
            if(_zz_357[62]) begin
              cntLkRespRmt_62 <= 6'h0;
            end
            if(_zz_357[63]) begin
              cntLkRespRmt_63 <= 6'h0;
            end
            if(_zz_358[0]) begin
              cntLkHoldLoc_0 <= 6'h0;
            end
            if(_zz_358[1]) begin
              cntLkHoldLoc_1 <= 6'h0;
            end
            if(_zz_358[2]) begin
              cntLkHoldLoc_2 <= 6'h0;
            end
            if(_zz_358[3]) begin
              cntLkHoldLoc_3 <= 6'h0;
            end
            if(_zz_358[4]) begin
              cntLkHoldLoc_4 <= 6'h0;
            end
            if(_zz_358[5]) begin
              cntLkHoldLoc_5 <= 6'h0;
            end
            if(_zz_358[6]) begin
              cntLkHoldLoc_6 <= 6'h0;
            end
            if(_zz_358[7]) begin
              cntLkHoldLoc_7 <= 6'h0;
            end
            if(_zz_358[8]) begin
              cntLkHoldLoc_8 <= 6'h0;
            end
            if(_zz_358[9]) begin
              cntLkHoldLoc_9 <= 6'h0;
            end
            if(_zz_358[10]) begin
              cntLkHoldLoc_10 <= 6'h0;
            end
            if(_zz_358[11]) begin
              cntLkHoldLoc_11 <= 6'h0;
            end
            if(_zz_358[12]) begin
              cntLkHoldLoc_12 <= 6'h0;
            end
            if(_zz_358[13]) begin
              cntLkHoldLoc_13 <= 6'h0;
            end
            if(_zz_358[14]) begin
              cntLkHoldLoc_14 <= 6'h0;
            end
            if(_zz_358[15]) begin
              cntLkHoldLoc_15 <= 6'h0;
            end
            if(_zz_358[16]) begin
              cntLkHoldLoc_16 <= 6'h0;
            end
            if(_zz_358[17]) begin
              cntLkHoldLoc_17 <= 6'h0;
            end
            if(_zz_358[18]) begin
              cntLkHoldLoc_18 <= 6'h0;
            end
            if(_zz_358[19]) begin
              cntLkHoldLoc_19 <= 6'h0;
            end
            if(_zz_358[20]) begin
              cntLkHoldLoc_20 <= 6'h0;
            end
            if(_zz_358[21]) begin
              cntLkHoldLoc_21 <= 6'h0;
            end
            if(_zz_358[22]) begin
              cntLkHoldLoc_22 <= 6'h0;
            end
            if(_zz_358[23]) begin
              cntLkHoldLoc_23 <= 6'h0;
            end
            if(_zz_358[24]) begin
              cntLkHoldLoc_24 <= 6'h0;
            end
            if(_zz_358[25]) begin
              cntLkHoldLoc_25 <= 6'h0;
            end
            if(_zz_358[26]) begin
              cntLkHoldLoc_26 <= 6'h0;
            end
            if(_zz_358[27]) begin
              cntLkHoldLoc_27 <= 6'h0;
            end
            if(_zz_358[28]) begin
              cntLkHoldLoc_28 <= 6'h0;
            end
            if(_zz_358[29]) begin
              cntLkHoldLoc_29 <= 6'h0;
            end
            if(_zz_358[30]) begin
              cntLkHoldLoc_30 <= 6'h0;
            end
            if(_zz_358[31]) begin
              cntLkHoldLoc_31 <= 6'h0;
            end
            if(_zz_358[32]) begin
              cntLkHoldLoc_32 <= 6'h0;
            end
            if(_zz_358[33]) begin
              cntLkHoldLoc_33 <= 6'h0;
            end
            if(_zz_358[34]) begin
              cntLkHoldLoc_34 <= 6'h0;
            end
            if(_zz_358[35]) begin
              cntLkHoldLoc_35 <= 6'h0;
            end
            if(_zz_358[36]) begin
              cntLkHoldLoc_36 <= 6'h0;
            end
            if(_zz_358[37]) begin
              cntLkHoldLoc_37 <= 6'h0;
            end
            if(_zz_358[38]) begin
              cntLkHoldLoc_38 <= 6'h0;
            end
            if(_zz_358[39]) begin
              cntLkHoldLoc_39 <= 6'h0;
            end
            if(_zz_358[40]) begin
              cntLkHoldLoc_40 <= 6'h0;
            end
            if(_zz_358[41]) begin
              cntLkHoldLoc_41 <= 6'h0;
            end
            if(_zz_358[42]) begin
              cntLkHoldLoc_42 <= 6'h0;
            end
            if(_zz_358[43]) begin
              cntLkHoldLoc_43 <= 6'h0;
            end
            if(_zz_358[44]) begin
              cntLkHoldLoc_44 <= 6'h0;
            end
            if(_zz_358[45]) begin
              cntLkHoldLoc_45 <= 6'h0;
            end
            if(_zz_358[46]) begin
              cntLkHoldLoc_46 <= 6'h0;
            end
            if(_zz_358[47]) begin
              cntLkHoldLoc_47 <= 6'h0;
            end
            if(_zz_358[48]) begin
              cntLkHoldLoc_48 <= 6'h0;
            end
            if(_zz_358[49]) begin
              cntLkHoldLoc_49 <= 6'h0;
            end
            if(_zz_358[50]) begin
              cntLkHoldLoc_50 <= 6'h0;
            end
            if(_zz_358[51]) begin
              cntLkHoldLoc_51 <= 6'h0;
            end
            if(_zz_358[52]) begin
              cntLkHoldLoc_52 <= 6'h0;
            end
            if(_zz_358[53]) begin
              cntLkHoldLoc_53 <= 6'h0;
            end
            if(_zz_358[54]) begin
              cntLkHoldLoc_54 <= 6'h0;
            end
            if(_zz_358[55]) begin
              cntLkHoldLoc_55 <= 6'h0;
            end
            if(_zz_358[56]) begin
              cntLkHoldLoc_56 <= 6'h0;
            end
            if(_zz_358[57]) begin
              cntLkHoldLoc_57 <= 6'h0;
            end
            if(_zz_358[58]) begin
              cntLkHoldLoc_58 <= 6'h0;
            end
            if(_zz_358[59]) begin
              cntLkHoldLoc_59 <= 6'h0;
            end
            if(_zz_358[60]) begin
              cntLkHoldLoc_60 <= 6'h0;
            end
            if(_zz_358[61]) begin
              cntLkHoldLoc_61 <= 6'h0;
            end
            if(_zz_358[62]) begin
              cntLkHoldLoc_62 <= 6'h0;
            end
            if(_zz_358[63]) begin
              cntLkHoldLoc_63 <= 6'h0;
            end
            if(_zz_359[0]) begin
              cntLkHoldRmt_0 <= 6'h0;
            end
            if(_zz_359[1]) begin
              cntLkHoldRmt_1 <= 6'h0;
            end
            if(_zz_359[2]) begin
              cntLkHoldRmt_2 <= 6'h0;
            end
            if(_zz_359[3]) begin
              cntLkHoldRmt_3 <= 6'h0;
            end
            if(_zz_359[4]) begin
              cntLkHoldRmt_4 <= 6'h0;
            end
            if(_zz_359[5]) begin
              cntLkHoldRmt_5 <= 6'h0;
            end
            if(_zz_359[6]) begin
              cntLkHoldRmt_6 <= 6'h0;
            end
            if(_zz_359[7]) begin
              cntLkHoldRmt_7 <= 6'h0;
            end
            if(_zz_359[8]) begin
              cntLkHoldRmt_8 <= 6'h0;
            end
            if(_zz_359[9]) begin
              cntLkHoldRmt_9 <= 6'h0;
            end
            if(_zz_359[10]) begin
              cntLkHoldRmt_10 <= 6'h0;
            end
            if(_zz_359[11]) begin
              cntLkHoldRmt_11 <= 6'h0;
            end
            if(_zz_359[12]) begin
              cntLkHoldRmt_12 <= 6'h0;
            end
            if(_zz_359[13]) begin
              cntLkHoldRmt_13 <= 6'h0;
            end
            if(_zz_359[14]) begin
              cntLkHoldRmt_14 <= 6'h0;
            end
            if(_zz_359[15]) begin
              cntLkHoldRmt_15 <= 6'h0;
            end
            if(_zz_359[16]) begin
              cntLkHoldRmt_16 <= 6'h0;
            end
            if(_zz_359[17]) begin
              cntLkHoldRmt_17 <= 6'h0;
            end
            if(_zz_359[18]) begin
              cntLkHoldRmt_18 <= 6'h0;
            end
            if(_zz_359[19]) begin
              cntLkHoldRmt_19 <= 6'h0;
            end
            if(_zz_359[20]) begin
              cntLkHoldRmt_20 <= 6'h0;
            end
            if(_zz_359[21]) begin
              cntLkHoldRmt_21 <= 6'h0;
            end
            if(_zz_359[22]) begin
              cntLkHoldRmt_22 <= 6'h0;
            end
            if(_zz_359[23]) begin
              cntLkHoldRmt_23 <= 6'h0;
            end
            if(_zz_359[24]) begin
              cntLkHoldRmt_24 <= 6'h0;
            end
            if(_zz_359[25]) begin
              cntLkHoldRmt_25 <= 6'h0;
            end
            if(_zz_359[26]) begin
              cntLkHoldRmt_26 <= 6'h0;
            end
            if(_zz_359[27]) begin
              cntLkHoldRmt_27 <= 6'h0;
            end
            if(_zz_359[28]) begin
              cntLkHoldRmt_28 <= 6'h0;
            end
            if(_zz_359[29]) begin
              cntLkHoldRmt_29 <= 6'h0;
            end
            if(_zz_359[30]) begin
              cntLkHoldRmt_30 <= 6'h0;
            end
            if(_zz_359[31]) begin
              cntLkHoldRmt_31 <= 6'h0;
            end
            if(_zz_359[32]) begin
              cntLkHoldRmt_32 <= 6'h0;
            end
            if(_zz_359[33]) begin
              cntLkHoldRmt_33 <= 6'h0;
            end
            if(_zz_359[34]) begin
              cntLkHoldRmt_34 <= 6'h0;
            end
            if(_zz_359[35]) begin
              cntLkHoldRmt_35 <= 6'h0;
            end
            if(_zz_359[36]) begin
              cntLkHoldRmt_36 <= 6'h0;
            end
            if(_zz_359[37]) begin
              cntLkHoldRmt_37 <= 6'h0;
            end
            if(_zz_359[38]) begin
              cntLkHoldRmt_38 <= 6'h0;
            end
            if(_zz_359[39]) begin
              cntLkHoldRmt_39 <= 6'h0;
            end
            if(_zz_359[40]) begin
              cntLkHoldRmt_40 <= 6'h0;
            end
            if(_zz_359[41]) begin
              cntLkHoldRmt_41 <= 6'h0;
            end
            if(_zz_359[42]) begin
              cntLkHoldRmt_42 <= 6'h0;
            end
            if(_zz_359[43]) begin
              cntLkHoldRmt_43 <= 6'h0;
            end
            if(_zz_359[44]) begin
              cntLkHoldRmt_44 <= 6'h0;
            end
            if(_zz_359[45]) begin
              cntLkHoldRmt_45 <= 6'h0;
            end
            if(_zz_359[46]) begin
              cntLkHoldRmt_46 <= 6'h0;
            end
            if(_zz_359[47]) begin
              cntLkHoldRmt_47 <= 6'h0;
            end
            if(_zz_359[48]) begin
              cntLkHoldRmt_48 <= 6'h0;
            end
            if(_zz_359[49]) begin
              cntLkHoldRmt_49 <= 6'h0;
            end
            if(_zz_359[50]) begin
              cntLkHoldRmt_50 <= 6'h0;
            end
            if(_zz_359[51]) begin
              cntLkHoldRmt_51 <= 6'h0;
            end
            if(_zz_359[52]) begin
              cntLkHoldRmt_52 <= 6'h0;
            end
            if(_zz_359[53]) begin
              cntLkHoldRmt_53 <= 6'h0;
            end
            if(_zz_359[54]) begin
              cntLkHoldRmt_54 <= 6'h0;
            end
            if(_zz_359[55]) begin
              cntLkHoldRmt_55 <= 6'h0;
            end
            if(_zz_359[56]) begin
              cntLkHoldRmt_56 <= 6'h0;
            end
            if(_zz_359[57]) begin
              cntLkHoldRmt_57 <= 6'h0;
            end
            if(_zz_359[58]) begin
              cntLkHoldRmt_58 <= 6'h0;
            end
            if(_zz_359[59]) begin
              cntLkHoldRmt_59 <= 6'h0;
            end
            if(_zz_359[60]) begin
              cntLkHoldRmt_60 <= 6'h0;
            end
            if(_zz_359[61]) begin
              cntLkHoldRmt_61 <= 6'h0;
            end
            if(_zz_359[62]) begin
              cntLkHoldRmt_62 <= 6'h0;
            end
            if(_zz_359[63]) begin
              cntLkHoldRmt_63 <= 6'h0;
            end
            if(_zz_360[0]) begin
              cntLkWaitLoc_0 <= 6'h0;
            end
            if(_zz_360[1]) begin
              cntLkWaitLoc_1 <= 6'h0;
            end
            if(_zz_360[2]) begin
              cntLkWaitLoc_2 <= 6'h0;
            end
            if(_zz_360[3]) begin
              cntLkWaitLoc_3 <= 6'h0;
            end
            if(_zz_360[4]) begin
              cntLkWaitLoc_4 <= 6'h0;
            end
            if(_zz_360[5]) begin
              cntLkWaitLoc_5 <= 6'h0;
            end
            if(_zz_360[6]) begin
              cntLkWaitLoc_6 <= 6'h0;
            end
            if(_zz_360[7]) begin
              cntLkWaitLoc_7 <= 6'h0;
            end
            if(_zz_360[8]) begin
              cntLkWaitLoc_8 <= 6'h0;
            end
            if(_zz_360[9]) begin
              cntLkWaitLoc_9 <= 6'h0;
            end
            if(_zz_360[10]) begin
              cntLkWaitLoc_10 <= 6'h0;
            end
            if(_zz_360[11]) begin
              cntLkWaitLoc_11 <= 6'h0;
            end
            if(_zz_360[12]) begin
              cntLkWaitLoc_12 <= 6'h0;
            end
            if(_zz_360[13]) begin
              cntLkWaitLoc_13 <= 6'h0;
            end
            if(_zz_360[14]) begin
              cntLkWaitLoc_14 <= 6'h0;
            end
            if(_zz_360[15]) begin
              cntLkWaitLoc_15 <= 6'h0;
            end
            if(_zz_360[16]) begin
              cntLkWaitLoc_16 <= 6'h0;
            end
            if(_zz_360[17]) begin
              cntLkWaitLoc_17 <= 6'h0;
            end
            if(_zz_360[18]) begin
              cntLkWaitLoc_18 <= 6'h0;
            end
            if(_zz_360[19]) begin
              cntLkWaitLoc_19 <= 6'h0;
            end
            if(_zz_360[20]) begin
              cntLkWaitLoc_20 <= 6'h0;
            end
            if(_zz_360[21]) begin
              cntLkWaitLoc_21 <= 6'h0;
            end
            if(_zz_360[22]) begin
              cntLkWaitLoc_22 <= 6'h0;
            end
            if(_zz_360[23]) begin
              cntLkWaitLoc_23 <= 6'h0;
            end
            if(_zz_360[24]) begin
              cntLkWaitLoc_24 <= 6'h0;
            end
            if(_zz_360[25]) begin
              cntLkWaitLoc_25 <= 6'h0;
            end
            if(_zz_360[26]) begin
              cntLkWaitLoc_26 <= 6'h0;
            end
            if(_zz_360[27]) begin
              cntLkWaitLoc_27 <= 6'h0;
            end
            if(_zz_360[28]) begin
              cntLkWaitLoc_28 <= 6'h0;
            end
            if(_zz_360[29]) begin
              cntLkWaitLoc_29 <= 6'h0;
            end
            if(_zz_360[30]) begin
              cntLkWaitLoc_30 <= 6'h0;
            end
            if(_zz_360[31]) begin
              cntLkWaitLoc_31 <= 6'h0;
            end
            if(_zz_360[32]) begin
              cntLkWaitLoc_32 <= 6'h0;
            end
            if(_zz_360[33]) begin
              cntLkWaitLoc_33 <= 6'h0;
            end
            if(_zz_360[34]) begin
              cntLkWaitLoc_34 <= 6'h0;
            end
            if(_zz_360[35]) begin
              cntLkWaitLoc_35 <= 6'h0;
            end
            if(_zz_360[36]) begin
              cntLkWaitLoc_36 <= 6'h0;
            end
            if(_zz_360[37]) begin
              cntLkWaitLoc_37 <= 6'h0;
            end
            if(_zz_360[38]) begin
              cntLkWaitLoc_38 <= 6'h0;
            end
            if(_zz_360[39]) begin
              cntLkWaitLoc_39 <= 6'h0;
            end
            if(_zz_360[40]) begin
              cntLkWaitLoc_40 <= 6'h0;
            end
            if(_zz_360[41]) begin
              cntLkWaitLoc_41 <= 6'h0;
            end
            if(_zz_360[42]) begin
              cntLkWaitLoc_42 <= 6'h0;
            end
            if(_zz_360[43]) begin
              cntLkWaitLoc_43 <= 6'h0;
            end
            if(_zz_360[44]) begin
              cntLkWaitLoc_44 <= 6'h0;
            end
            if(_zz_360[45]) begin
              cntLkWaitLoc_45 <= 6'h0;
            end
            if(_zz_360[46]) begin
              cntLkWaitLoc_46 <= 6'h0;
            end
            if(_zz_360[47]) begin
              cntLkWaitLoc_47 <= 6'h0;
            end
            if(_zz_360[48]) begin
              cntLkWaitLoc_48 <= 6'h0;
            end
            if(_zz_360[49]) begin
              cntLkWaitLoc_49 <= 6'h0;
            end
            if(_zz_360[50]) begin
              cntLkWaitLoc_50 <= 6'h0;
            end
            if(_zz_360[51]) begin
              cntLkWaitLoc_51 <= 6'h0;
            end
            if(_zz_360[52]) begin
              cntLkWaitLoc_52 <= 6'h0;
            end
            if(_zz_360[53]) begin
              cntLkWaitLoc_53 <= 6'h0;
            end
            if(_zz_360[54]) begin
              cntLkWaitLoc_54 <= 6'h0;
            end
            if(_zz_360[55]) begin
              cntLkWaitLoc_55 <= 6'h0;
            end
            if(_zz_360[56]) begin
              cntLkWaitLoc_56 <= 6'h0;
            end
            if(_zz_360[57]) begin
              cntLkWaitLoc_57 <= 6'h0;
            end
            if(_zz_360[58]) begin
              cntLkWaitLoc_58 <= 6'h0;
            end
            if(_zz_360[59]) begin
              cntLkWaitLoc_59 <= 6'h0;
            end
            if(_zz_360[60]) begin
              cntLkWaitLoc_60 <= 6'h0;
            end
            if(_zz_360[61]) begin
              cntLkWaitLoc_61 <= 6'h0;
            end
            if(_zz_360[62]) begin
              cntLkWaitLoc_62 <= 6'h0;
            end
            if(_zz_360[63]) begin
              cntLkWaitLoc_63 <= 6'h0;
            end
            if(_zz_361[0]) begin
              cntLkWaitRmt_0 <= 6'h0;
            end
            if(_zz_361[1]) begin
              cntLkWaitRmt_1 <= 6'h0;
            end
            if(_zz_361[2]) begin
              cntLkWaitRmt_2 <= 6'h0;
            end
            if(_zz_361[3]) begin
              cntLkWaitRmt_3 <= 6'h0;
            end
            if(_zz_361[4]) begin
              cntLkWaitRmt_4 <= 6'h0;
            end
            if(_zz_361[5]) begin
              cntLkWaitRmt_5 <= 6'h0;
            end
            if(_zz_361[6]) begin
              cntLkWaitRmt_6 <= 6'h0;
            end
            if(_zz_361[7]) begin
              cntLkWaitRmt_7 <= 6'h0;
            end
            if(_zz_361[8]) begin
              cntLkWaitRmt_8 <= 6'h0;
            end
            if(_zz_361[9]) begin
              cntLkWaitRmt_9 <= 6'h0;
            end
            if(_zz_361[10]) begin
              cntLkWaitRmt_10 <= 6'h0;
            end
            if(_zz_361[11]) begin
              cntLkWaitRmt_11 <= 6'h0;
            end
            if(_zz_361[12]) begin
              cntLkWaitRmt_12 <= 6'h0;
            end
            if(_zz_361[13]) begin
              cntLkWaitRmt_13 <= 6'h0;
            end
            if(_zz_361[14]) begin
              cntLkWaitRmt_14 <= 6'h0;
            end
            if(_zz_361[15]) begin
              cntLkWaitRmt_15 <= 6'h0;
            end
            if(_zz_361[16]) begin
              cntLkWaitRmt_16 <= 6'h0;
            end
            if(_zz_361[17]) begin
              cntLkWaitRmt_17 <= 6'h0;
            end
            if(_zz_361[18]) begin
              cntLkWaitRmt_18 <= 6'h0;
            end
            if(_zz_361[19]) begin
              cntLkWaitRmt_19 <= 6'h0;
            end
            if(_zz_361[20]) begin
              cntLkWaitRmt_20 <= 6'h0;
            end
            if(_zz_361[21]) begin
              cntLkWaitRmt_21 <= 6'h0;
            end
            if(_zz_361[22]) begin
              cntLkWaitRmt_22 <= 6'h0;
            end
            if(_zz_361[23]) begin
              cntLkWaitRmt_23 <= 6'h0;
            end
            if(_zz_361[24]) begin
              cntLkWaitRmt_24 <= 6'h0;
            end
            if(_zz_361[25]) begin
              cntLkWaitRmt_25 <= 6'h0;
            end
            if(_zz_361[26]) begin
              cntLkWaitRmt_26 <= 6'h0;
            end
            if(_zz_361[27]) begin
              cntLkWaitRmt_27 <= 6'h0;
            end
            if(_zz_361[28]) begin
              cntLkWaitRmt_28 <= 6'h0;
            end
            if(_zz_361[29]) begin
              cntLkWaitRmt_29 <= 6'h0;
            end
            if(_zz_361[30]) begin
              cntLkWaitRmt_30 <= 6'h0;
            end
            if(_zz_361[31]) begin
              cntLkWaitRmt_31 <= 6'h0;
            end
            if(_zz_361[32]) begin
              cntLkWaitRmt_32 <= 6'h0;
            end
            if(_zz_361[33]) begin
              cntLkWaitRmt_33 <= 6'h0;
            end
            if(_zz_361[34]) begin
              cntLkWaitRmt_34 <= 6'h0;
            end
            if(_zz_361[35]) begin
              cntLkWaitRmt_35 <= 6'h0;
            end
            if(_zz_361[36]) begin
              cntLkWaitRmt_36 <= 6'h0;
            end
            if(_zz_361[37]) begin
              cntLkWaitRmt_37 <= 6'h0;
            end
            if(_zz_361[38]) begin
              cntLkWaitRmt_38 <= 6'h0;
            end
            if(_zz_361[39]) begin
              cntLkWaitRmt_39 <= 6'h0;
            end
            if(_zz_361[40]) begin
              cntLkWaitRmt_40 <= 6'h0;
            end
            if(_zz_361[41]) begin
              cntLkWaitRmt_41 <= 6'h0;
            end
            if(_zz_361[42]) begin
              cntLkWaitRmt_42 <= 6'h0;
            end
            if(_zz_361[43]) begin
              cntLkWaitRmt_43 <= 6'h0;
            end
            if(_zz_361[44]) begin
              cntLkWaitRmt_44 <= 6'h0;
            end
            if(_zz_361[45]) begin
              cntLkWaitRmt_45 <= 6'h0;
            end
            if(_zz_361[46]) begin
              cntLkWaitRmt_46 <= 6'h0;
            end
            if(_zz_361[47]) begin
              cntLkWaitRmt_47 <= 6'h0;
            end
            if(_zz_361[48]) begin
              cntLkWaitRmt_48 <= 6'h0;
            end
            if(_zz_361[49]) begin
              cntLkWaitRmt_49 <= 6'h0;
            end
            if(_zz_361[50]) begin
              cntLkWaitRmt_50 <= 6'h0;
            end
            if(_zz_361[51]) begin
              cntLkWaitRmt_51 <= 6'h0;
            end
            if(_zz_361[52]) begin
              cntLkWaitRmt_52 <= 6'h0;
            end
            if(_zz_361[53]) begin
              cntLkWaitRmt_53 <= 6'h0;
            end
            if(_zz_361[54]) begin
              cntLkWaitRmt_54 <= 6'h0;
            end
            if(_zz_361[55]) begin
              cntLkWaitRmt_55 <= 6'h0;
            end
            if(_zz_361[56]) begin
              cntLkWaitRmt_56 <= 6'h0;
            end
            if(_zz_361[57]) begin
              cntLkWaitRmt_57 <= 6'h0;
            end
            if(_zz_361[58]) begin
              cntLkWaitRmt_58 <= 6'h0;
            end
            if(_zz_361[59]) begin
              cntLkWaitRmt_59 <= 6'h0;
            end
            if(_zz_361[60]) begin
              cntLkWaitRmt_60 <= 6'h0;
            end
            if(_zz_361[61]) begin
              cntLkWaitRmt_61 <= 6'h0;
            end
            if(_zz_361[62]) begin
              cntLkWaitRmt_62 <= 6'h0;
            end
            if(_zz_361[63]) begin
              cntLkWaitRmt_63 <= 6'h0;
            end
            if(_zz_362[0]) begin
              cntLkReqWrLoc_0 <= 6'h0;
            end
            if(_zz_362[1]) begin
              cntLkReqWrLoc_1 <= 6'h0;
            end
            if(_zz_362[2]) begin
              cntLkReqWrLoc_2 <= 6'h0;
            end
            if(_zz_362[3]) begin
              cntLkReqWrLoc_3 <= 6'h0;
            end
            if(_zz_362[4]) begin
              cntLkReqWrLoc_4 <= 6'h0;
            end
            if(_zz_362[5]) begin
              cntLkReqWrLoc_5 <= 6'h0;
            end
            if(_zz_362[6]) begin
              cntLkReqWrLoc_6 <= 6'h0;
            end
            if(_zz_362[7]) begin
              cntLkReqWrLoc_7 <= 6'h0;
            end
            if(_zz_362[8]) begin
              cntLkReqWrLoc_8 <= 6'h0;
            end
            if(_zz_362[9]) begin
              cntLkReqWrLoc_9 <= 6'h0;
            end
            if(_zz_362[10]) begin
              cntLkReqWrLoc_10 <= 6'h0;
            end
            if(_zz_362[11]) begin
              cntLkReqWrLoc_11 <= 6'h0;
            end
            if(_zz_362[12]) begin
              cntLkReqWrLoc_12 <= 6'h0;
            end
            if(_zz_362[13]) begin
              cntLkReqWrLoc_13 <= 6'h0;
            end
            if(_zz_362[14]) begin
              cntLkReqWrLoc_14 <= 6'h0;
            end
            if(_zz_362[15]) begin
              cntLkReqWrLoc_15 <= 6'h0;
            end
            if(_zz_362[16]) begin
              cntLkReqWrLoc_16 <= 6'h0;
            end
            if(_zz_362[17]) begin
              cntLkReqWrLoc_17 <= 6'h0;
            end
            if(_zz_362[18]) begin
              cntLkReqWrLoc_18 <= 6'h0;
            end
            if(_zz_362[19]) begin
              cntLkReqWrLoc_19 <= 6'h0;
            end
            if(_zz_362[20]) begin
              cntLkReqWrLoc_20 <= 6'h0;
            end
            if(_zz_362[21]) begin
              cntLkReqWrLoc_21 <= 6'h0;
            end
            if(_zz_362[22]) begin
              cntLkReqWrLoc_22 <= 6'h0;
            end
            if(_zz_362[23]) begin
              cntLkReqWrLoc_23 <= 6'h0;
            end
            if(_zz_362[24]) begin
              cntLkReqWrLoc_24 <= 6'h0;
            end
            if(_zz_362[25]) begin
              cntLkReqWrLoc_25 <= 6'h0;
            end
            if(_zz_362[26]) begin
              cntLkReqWrLoc_26 <= 6'h0;
            end
            if(_zz_362[27]) begin
              cntLkReqWrLoc_27 <= 6'h0;
            end
            if(_zz_362[28]) begin
              cntLkReqWrLoc_28 <= 6'h0;
            end
            if(_zz_362[29]) begin
              cntLkReqWrLoc_29 <= 6'h0;
            end
            if(_zz_362[30]) begin
              cntLkReqWrLoc_30 <= 6'h0;
            end
            if(_zz_362[31]) begin
              cntLkReqWrLoc_31 <= 6'h0;
            end
            if(_zz_362[32]) begin
              cntLkReqWrLoc_32 <= 6'h0;
            end
            if(_zz_362[33]) begin
              cntLkReqWrLoc_33 <= 6'h0;
            end
            if(_zz_362[34]) begin
              cntLkReqWrLoc_34 <= 6'h0;
            end
            if(_zz_362[35]) begin
              cntLkReqWrLoc_35 <= 6'h0;
            end
            if(_zz_362[36]) begin
              cntLkReqWrLoc_36 <= 6'h0;
            end
            if(_zz_362[37]) begin
              cntLkReqWrLoc_37 <= 6'h0;
            end
            if(_zz_362[38]) begin
              cntLkReqWrLoc_38 <= 6'h0;
            end
            if(_zz_362[39]) begin
              cntLkReqWrLoc_39 <= 6'h0;
            end
            if(_zz_362[40]) begin
              cntLkReqWrLoc_40 <= 6'h0;
            end
            if(_zz_362[41]) begin
              cntLkReqWrLoc_41 <= 6'h0;
            end
            if(_zz_362[42]) begin
              cntLkReqWrLoc_42 <= 6'h0;
            end
            if(_zz_362[43]) begin
              cntLkReqWrLoc_43 <= 6'h0;
            end
            if(_zz_362[44]) begin
              cntLkReqWrLoc_44 <= 6'h0;
            end
            if(_zz_362[45]) begin
              cntLkReqWrLoc_45 <= 6'h0;
            end
            if(_zz_362[46]) begin
              cntLkReqWrLoc_46 <= 6'h0;
            end
            if(_zz_362[47]) begin
              cntLkReqWrLoc_47 <= 6'h0;
            end
            if(_zz_362[48]) begin
              cntLkReqWrLoc_48 <= 6'h0;
            end
            if(_zz_362[49]) begin
              cntLkReqWrLoc_49 <= 6'h0;
            end
            if(_zz_362[50]) begin
              cntLkReqWrLoc_50 <= 6'h0;
            end
            if(_zz_362[51]) begin
              cntLkReqWrLoc_51 <= 6'h0;
            end
            if(_zz_362[52]) begin
              cntLkReqWrLoc_52 <= 6'h0;
            end
            if(_zz_362[53]) begin
              cntLkReqWrLoc_53 <= 6'h0;
            end
            if(_zz_362[54]) begin
              cntLkReqWrLoc_54 <= 6'h0;
            end
            if(_zz_362[55]) begin
              cntLkReqWrLoc_55 <= 6'h0;
            end
            if(_zz_362[56]) begin
              cntLkReqWrLoc_56 <= 6'h0;
            end
            if(_zz_362[57]) begin
              cntLkReqWrLoc_57 <= 6'h0;
            end
            if(_zz_362[58]) begin
              cntLkReqWrLoc_58 <= 6'h0;
            end
            if(_zz_362[59]) begin
              cntLkReqWrLoc_59 <= 6'h0;
            end
            if(_zz_362[60]) begin
              cntLkReqWrLoc_60 <= 6'h0;
            end
            if(_zz_362[61]) begin
              cntLkReqWrLoc_61 <= 6'h0;
            end
            if(_zz_362[62]) begin
              cntLkReqWrLoc_62 <= 6'h0;
            end
            if(_zz_362[63]) begin
              cntLkReqWrLoc_63 <= 6'h0;
            end
            if(_zz_363[0]) begin
              cntLkReqWrRmt_0 <= 6'h0;
            end
            if(_zz_363[1]) begin
              cntLkReqWrRmt_1 <= 6'h0;
            end
            if(_zz_363[2]) begin
              cntLkReqWrRmt_2 <= 6'h0;
            end
            if(_zz_363[3]) begin
              cntLkReqWrRmt_3 <= 6'h0;
            end
            if(_zz_363[4]) begin
              cntLkReqWrRmt_4 <= 6'h0;
            end
            if(_zz_363[5]) begin
              cntLkReqWrRmt_5 <= 6'h0;
            end
            if(_zz_363[6]) begin
              cntLkReqWrRmt_6 <= 6'h0;
            end
            if(_zz_363[7]) begin
              cntLkReqWrRmt_7 <= 6'h0;
            end
            if(_zz_363[8]) begin
              cntLkReqWrRmt_8 <= 6'h0;
            end
            if(_zz_363[9]) begin
              cntLkReqWrRmt_9 <= 6'h0;
            end
            if(_zz_363[10]) begin
              cntLkReqWrRmt_10 <= 6'h0;
            end
            if(_zz_363[11]) begin
              cntLkReqWrRmt_11 <= 6'h0;
            end
            if(_zz_363[12]) begin
              cntLkReqWrRmt_12 <= 6'h0;
            end
            if(_zz_363[13]) begin
              cntLkReqWrRmt_13 <= 6'h0;
            end
            if(_zz_363[14]) begin
              cntLkReqWrRmt_14 <= 6'h0;
            end
            if(_zz_363[15]) begin
              cntLkReqWrRmt_15 <= 6'h0;
            end
            if(_zz_363[16]) begin
              cntLkReqWrRmt_16 <= 6'h0;
            end
            if(_zz_363[17]) begin
              cntLkReqWrRmt_17 <= 6'h0;
            end
            if(_zz_363[18]) begin
              cntLkReqWrRmt_18 <= 6'h0;
            end
            if(_zz_363[19]) begin
              cntLkReqWrRmt_19 <= 6'h0;
            end
            if(_zz_363[20]) begin
              cntLkReqWrRmt_20 <= 6'h0;
            end
            if(_zz_363[21]) begin
              cntLkReqWrRmt_21 <= 6'h0;
            end
            if(_zz_363[22]) begin
              cntLkReqWrRmt_22 <= 6'h0;
            end
            if(_zz_363[23]) begin
              cntLkReqWrRmt_23 <= 6'h0;
            end
            if(_zz_363[24]) begin
              cntLkReqWrRmt_24 <= 6'h0;
            end
            if(_zz_363[25]) begin
              cntLkReqWrRmt_25 <= 6'h0;
            end
            if(_zz_363[26]) begin
              cntLkReqWrRmt_26 <= 6'h0;
            end
            if(_zz_363[27]) begin
              cntLkReqWrRmt_27 <= 6'h0;
            end
            if(_zz_363[28]) begin
              cntLkReqWrRmt_28 <= 6'h0;
            end
            if(_zz_363[29]) begin
              cntLkReqWrRmt_29 <= 6'h0;
            end
            if(_zz_363[30]) begin
              cntLkReqWrRmt_30 <= 6'h0;
            end
            if(_zz_363[31]) begin
              cntLkReqWrRmt_31 <= 6'h0;
            end
            if(_zz_363[32]) begin
              cntLkReqWrRmt_32 <= 6'h0;
            end
            if(_zz_363[33]) begin
              cntLkReqWrRmt_33 <= 6'h0;
            end
            if(_zz_363[34]) begin
              cntLkReqWrRmt_34 <= 6'h0;
            end
            if(_zz_363[35]) begin
              cntLkReqWrRmt_35 <= 6'h0;
            end
            if(_zz_363[36]) begin
              cntLkReqWrRmt_36 <= 6'h0;
            end
            if(_zz_363[37]) begin
              cntLkReqWrRmt_37 <= 6'h0;
            end
            if(_zz_363[38]) begin
              cntLkReqWrRmt_38 <= 6'h0;
            end
            if(_zz_363[39]) begin
              cntLkReqWrRmt_39 <= 6'h0;
            end
            if(_zz_363[40]) begin
              cntLkReqWrRmt_40 <= 6'h0;
            end
            if(_zz_363[41]) begin
              cntLkReqWrRmt_41 <= 6'h0;
            end
            if(_zz_363[42]) begin
              cntLkReqWrRmt_42 <= 6'h0;
            end
            if(_zz_363[43]) begin
              cntLkReqWrRmt_43 <= 6'h0;
            end
            if(_zz_363[44]) begin
              cntLkReqWrRmt_44 <= 6'h0;
            end
            if(_zz_363[45]) begin
              cntLkReqWrRmt_45 <= 6'h0;
            end
            if(_zz_363[46]) begin
              cntLkReqWrRmt_46 <= 6'h0;
            end
            if(_zz_363[47]) begin
              cntLkReqWrRmt_47 <= 6'h0;
            end
            if(_zz_363[48]) begin
              cntLkReqWrRmt_48 <= 6'h0;
            end
            if(_zz_363[49]) begin
              cntLkReqWrRmt_49 <= 6'h0;
            end
            if(_zz_363[50]) begin
              cntLkReqWrRmt_50 <= 6'h0;
            end
            if(_zz_363[51]) begin
              cntLkReqWrRmt_51 <= 6'h0;
            end
            if(_zz_363[52]) begin
              cntLkReqWrRmt_52 <= 6'h0;
            end
            if(_zz_363[53]) begin
              cntLkReqWrRmt_53 <= 6'h0;
            end
            if(_zz_363[54]) begin
              cntLkReqWrRmt_54 <= 6'h0;
            end
            if(_zz_363[55]) begin
              cntLkReqWrRmt_55 <= 6'h0;
            end
            if(_zz_363[56]) begin
              cntLkReqWrRmt_56 <= 6'h0;
            end
            if(_zz_363[57]) begin
              cntLkReqWrRmt_57 <= 6'h0;
            end
            if(_zz_363[58]) begin
              cntLkReqWrRmt_58 <= 6'h0;
            end
            if(_zz_363[59]) begin
              cntLkReqWrRmt_59 <= 6'h0;
            end
            if(_zz_363[60]) begin
              cntLkReqWrRmt_60 <= 6'h0;
            end
            if(_zz_363[61]) begin
              cntLkReqWrRmt_61 <= 6'h0;
            end
            if(_zz_363[62]) begin
              cntLkReqWrRmt_62 <= 6'h0;
            end
            if(_zz_363[63]) begin
              cntLkReqWrRmt_63 <= 6'h0;
            end
            if(_zz_364[0]) begin
              cntLkHoldWrLoc_0 <= 6'h0;
            end
            if(_zz_364[1]) begin
              cntLkHoldWrLoc_1 <= 6'h0;
            end
            if(_zz_364[2]) begin
              cntLkHoldWrLoc_2 <= 6'h0;
            end
            if(_zz_364[3]) begin
              cntLkHoldWrLoc_3 <= 6'h0;
            end
            if(_zz_364[4]) begin
              cntLkHoldWrLoc_4 <= 6'h0;
            end
            if(_zz_364[5]) begin
              cntLkHoldWrLoc_5 <= 6'h0;
            end
            if(_zz_364[6]) begin
              cntLkHoldWrLoc_6 <= 6'h0;
            end
            if(_zz_364[7]) begin
              cntLkHoldWrLoc_7 <= 6'h0;
            end
            if(_zz_364[8]) begin
              cntLkHoldWrLoc_8 <= 6'h0;
            end
            if(_zz_364[9]) begin
              cntLkHoldWrLoc_9 <= 6'h0;
            end
            if(_zz_364[10]) begin
              cntLkHoldWrLoc_10 <= 6'h0;
            end
            if(_zz_364[11]) begin
              cntLkHoldWrLoc_11 <= 6'h0;
            end
            if(_zz_364[12]) begin
              cntLkHoldWrLoc_12 <= 6'h0;
            end
            if(_zz_364[13]) begin
              cntLkHoldWrLoc_13 <= 6'h0;
            end
            if(_zz_364[14]) begin
              cntLkHoldWrLoc_14 <= 6'h0;
            end
            if(_zz_364[15]) begin
              cntLkHoldWrLoc_15 <= 6'h0;
            end
            if(_zz_364[16]) begin
              cntLkHoldWrLoc_16 <= 6'h0;
            end
            if(_zz_364[17]) begin
              cntLkHoldWrLoc_17 <= 6'h0;
            end
            if(_zz_364[18]) begin
              cntLkHoldWrLoc_18 <= 6'h0;
            end
            if(_zz_364[19]) begin
              cntLkHoldWrLoc_19 <= 6'h0;
            end
            if(_zz_364[20]) begin
              cntLkHoldWrLoc_20 <= 6'h0;
            end
            if(_zz_364[21]) begin
              cntLkHoldWrLoc_21 <= 6'h0;
            end
            if(_zz_364[22]) begin
              cntLkHoldWrLoc_22 <= 6'h0;
            end
            if(_zz_364[23]) begin
              cntLkHoldWrLoc_23 <= 6'h0;
            end
            if(_zz_364[24]) begin
              cntLkHoldWrLoc_24 <= 6'h0;
            end
            if(_zz_364[25]) begin
              cntLkHoldWrLoc_25 <= 6'h0;
            end
            if(_zz_364[26]) begin
              cntLkHoldWrLoc_26 <= 6'h0;
            end
            if(_zz_364[27]) begin
              cntLkHoldWrLoc_27 <= 6'h0;
            end
            if(_zz_364[28]) begin
              cntLkHoldWrLoc_28 <= 6'h0;
            end
            if(_zz_364[29]) begin
              cntLkHoldWrLoc_29 <= 6'h0;
            end
            if(_zz_364[30]) begin
              cntLkHoldWrLoc_30 <= 6'h0;
            end
            if(_zz_364[31]) begin
              cntLkHoldWrLoc_31 <= 6'h0;
            end
            if(_zz_364[32]) begin
              cntLkHoldWrLoc_32 <= 6'h0;
            end
            if(_zz_364[33]) begin
              cntLkHoldWrLoc_33 <= 6'h0;
            end
            if(_zz_364[34]) begin
              cntLkHoldWrLoc_34 <= 6'h0;
            end
            if(_zz_364[35]) begin
              cntLkHoldWrLoc_35 <= 6'h0;
            end
            if(_zz_364[36]) begin
              cntLkHoldWrLoc_36 <= 6'h0;
            end
            if(_zz_364[37]) begin
              cntLkHoldWrLoc_37 <= 6'h0;
            end
            if(_zz_364[38]) begin
              cntLkHoldWrLoc_38 <= 6'h0;
            end
            if(_zz_364[39]) begin
              cntLkHoldWrLoc_39 <= 6'h0;
            end
            if(_zz_364[40]) begin
              cntLkHoldWrLoc_40 <= 6'h0;
            end
            if(_zz_364[41]) begin
              cntLkHoldWrLoc_41 <= 6'h0;
            end
            if(_zz_364[42]) begin
              cntLkHoldWrLoc_42 <= 6'h0;
            end
            if(_zz_364[43]) begin
              cntLkHoldWrLoc_43 <= 6'h0;
            end
            if(_zz_364[44]) begin
              cntLkHoldWrLoc_44 <= 6'h0;
            end
            if(_zz_364[45]) begin
              cntLkHoldWrLoc_45 <= 6'h0;
            end
            if(_zz_364[46]) begin
              cntLkHoldWrLoc_46 <= 6'h0;
            end
            if(_zz_364[47]) begin
              cntLkHoldWrLoc_47 <= 6'h0;
            end
            if(_zz_364[48]) begin
              cntLkHoldWrLoc_48 <= 6'h0;
            end
            if(_zz_364[49]) begin
              cntLkHoldWrLoc_49 <= 6'h0;
            end
            if(_zz_364[50]) begin
              cntLkHoldWrLoc_50 <= 6'h0;
            end
            if(_zz_364[51]) begin
              cntLkHoldWrLoc_51 <= 6'h0;
            end
            if(_zz_364[52]) begin
              cntLkHoldWrLoc_52 <= 6'h0;
            end
            if(_zz_364[53]) begin
              cntLkHoldWrLoc_53 <= 6'h0;
            end
            if(_zz_364[54]) begin
              cntLkHoldWrLoc_54 <= 6'h0;
            end
            if(_zz_364[55]) begin
              cntLkHoldWrLoc_55 <= 6'h0;
            end
            if(_zz_364[56]) begin
              cntLkHoldWrLoc_56 <= 6'h0;
            end
            if(_zz_364[57]) begin
              cntLkHoldWrLoc_57 <= 6'h0;
            end
            if(_zz_364[58]) begin
              cntLkHoldWrLoc_58 <= 6'h0;
            end
            if(_zz_364[59]) begin
              cntLkHoldWrLoc_59 <= 6'h0;
            end
            if(_zz_364[60]) begin
              cntLkHoldWrLoc_60 <= 6'h0;
            end
            if(_zz_364[61]) begin
              cntLkHoldWrLoc_61 <= 6'h0;
            end
            if(_zz_364[62]) begin
              cntLkHoldWrLoc_62 <= 6'h0;
            end
            if(_zz_364[63]) begin
              cntLkHoldWrLoc_63 <= 6'h0;
            end
            if(_zz_365[0]) begin
              cntLkHoldWrRmt_0 <= 6'h0;
            end
            if(_zz_365[1]) begin
              cntLkHoldWrRmt_1 <= 6'h0;
            end
            if(_zz_365[2]) begin
              cntLkHoldWrRmt_2 <= 6'h0;
            end
            if(_zz_365[3]) begin
              cntLkHoldWrRmt_3 <= 6'h0;
            end
            if(_zz_365[4]) begin
              cntLkHoldWrRmt_4 <= 6'h0;
            end
            if(_zz_365[5]) begin
              cntLkHoldWrRmt_5 <= 6'h0;
            end
            if(_zz_365[6]) begin
              cntLkHoldWrRmt_6 <= 6'h0;
            end
            if(_zz_365[7]) begin
              cntLkHoldWrRmt_7 <= 6'h0;
            end
            if(_zz_365[8]) begin
              cntLkHoldWrRmt_8 <= 6'h0;
            end
            if(_zz_365[9]) begin
              cntLkHoldWrRmt_9 <= 6'h0;
            end
            if(_zz_365[10]) begin
              cntLkHoldWrRmt_10 <= 6'h0;
            end
            if(_zz_365[11]) begin
              cntLkHoldWrRmt_11 <= 6'h0;
            end
            if(_zz_365[12]) begin
              cntLkHoldWrRmt_12 <= 6'h0;
            end
            if(_zz_365[13]) begin
              cntLkHoldWrRmt_13 <= 6'h0;
            end
            if(_zz_365[14]) begin
              cntLkHoldWrRmt_14 <= 6'h0;
            end
            if(_zz_365[15]) begin
              cntLkHoldWrRmt_15 <= 6'h0;
            end
            if(_zz_365[16]) begin
              cntLkHoldWrRmt_16 <= 6'h0;
            end
            if(_zz_365[17]) begin
              cntLkHoldWrRmt_17 <= 6'h0;
            end
            if(_zz_365[18]) begin
              cntLkHoldWrRmt_18 <= 6'h0;
            end
            if(_zz_365[19]) begin
              cntLkHoldWrRmt_19 <= 6'h0;
            end
            if(_zz_365[20]) begin
              cntLkHoldWrRmt_20 <= 6'h0;
            end
            if(_zz_365[21]) begin
              cntLkHoldWrRmt_21 <= 6'h0;
            end
            if(_zz_365[22]) begin
              cntLkHoldWrRmt_22 <= 6'h0;
            end
            if(_zz_365[23]) begin
              cntLkHoldWrRmt_23 <= 6'h0;
            end
            if(_zz_365[24]) begin
              cntLkHoldWrRmt_24 <= 6'h0;
            end
            if(_zz_365[25]) begin
              cntLkHoldWrRmt_25 <= 6'h0;
            end
            if(_zz_365[26]) begin
              cntLkHoldWrRmt_26 <= 6'h0;
            end
            if(_zz_365[27]) begin
              cntLkHoldWrRmt_27 <= 6'h0;
            end
            if(_zz_365[28]) begin
              cntLkHoldWrRmt_28 <= 6'h0;
            end
            if(_zz_365[29]) begin
              cntLkHoldWrRmt_29 <= 6'h0;
            end
            if(_zz_365[30]) begin
              cntLkHoldWrRmt_30 <= 6'h0;
            end
            if(_zz_365[31]) begin
              cntLkHoldWrRmt_31 <= 6'h0;
            end
            if(_zz_365[32]) begin
              cntLkHoldWrRmt_32 <= 6'h0;
            end
            if(_zz_365[33]) begin
              cntLkHoldWrRmt_33 <= 6'h0;
            end
            if(_zz_365[34]) begin
              cntLkHoldWrRmt_34 <= 6'h0;
            end
            if(_zz_365[35]) begin
              cntLkHoldWrRmt_35 <= 6'h0;
            end
            if(_zz_365[36]) begin
              cntLkHoldWrRmt_36 <= 6'h0;
            end
            if(_zz_365[37]) begin
              cntLkHoldWrRmt_37 <= 6'h0;
            end
            if(_zz_365[38]) begin
              cntLkHoldWrRmt_38 <= 6'h0;
            end
            if(_zz_365[39]) begin
              cntLkHoldWrRmt_39 <= 6'h0;
            end
            if(_zz_365[40]) begin
              cntLkHoldWrRmt_40 <= 6'h0;
            end
            if(_zz_365[41]) begin
              cntLkHoldWrRmt_41 <= 6'h0;
            end
            if(_zz_365[42]) begin
              cntLkHoldWrRmt_42 <= 6'h0;
            end
            if(_zz_365[43]) begin
              cntLkHoldWrRmt_43 <= 6'h0;
            end
            if(_zz_365[44]) begin
              cntLkHoldWrRmt_44 <= 6'h0;
            end
            if(_zz_365[45]) begin
              cntLkHoldWrRmt_45 <= 6'h0;
            end
            if(_zz_365[46]) begin
              cntLkHoldWrRmt_46 <= 6'h0;
            end
            if(_zz_365[47]) begin
              cntLkHoldWrRmt_47 <= 6'h0;
            end
            if(_zz_365[48]) begin
              cntLkHoldWrRmt_48 <= 6'h0;
            end
            if(_zz_365[49]) begin
              cntLkHoldWrRmt_49 <= 6'h0;
            end
            if(_zz_365[50]) begin
              cntLkHoldWrRmt_50 <= 6'h0;
            end
            if(_zz_365[51]) begin
              cntLkHoldWrRmt_51 <= 6'h0;
            end
            if(_zz_365[52]) begin
              cntLkHoldWrRmt_52 <= 6'h0;
            end
            if(_zz_365[53]) begin
              cntLkHoldWrRmt_53 <= 6'h0;
            end
            if(_zz_365[54]) begin
              cntLkHoldWrRmt_54 <= 6'h0;
            end
            if(_zz_365[55]) begin
              cntLkHoldWrRmt_55 <= 6'h0;
            end
            if(_zz_365[56]) begin
              cntLkHoldWrRmt_56 <= 6'h0;
            end
            if(_zz_365[57]) begin
              cntLkHoldWrRmt_57 <= 6'h0;
            end
            if(_zz_365[58]) begin
              cntLkHoldWrRmt_58 <= 6'h0;
            end
            if(_zz_365[59]) begin
              cntLkHoldWrRmt_59 <= 6'h0;
            end
            if(_zz_365[60]) begin
              cntLkHoldWrRmt_60 <= 6'h0;
            end
            if(_zz_365[61]) begin
              cntLkHoldWrRmt_61 <= 6'h0;
            end
            if(_zz_365[62]) begin
              cntLkHoldWrRmt_62 <= 6'h0;
            end
            if(_zz_365[63]) begin
              cntLkHoldWrRmt_63 <= 6'h0;
            end
            if(_zz_366[0]) begin
              cntCmtReqLoc_0 <= 6'h0;
            end
            if(_zz_366[1]) begin
              cntCmtReqLoc_1 <= 6'h0;
            end
            if(_zz_366[2]) begin
              cntCmtReqLoc_2 <= 6'h0;
            end
            if(_zz_366[3]) begin
              cntCmtReqLoc_3 <= 6'h0;
            end
            if(_zz_366[4]) begin
              cntCmtReqLoc_4 <= 6'h0;
            end
            if(_zz_366[5]) begin
              cntCmtReqLoc_5 <= 6'h0;
            end
            if(_zz_366[6]) begin
              cntCmtReqLoc_6 <= 6'h0;
            end
            if(_zz_366[7]) begin
              cntCmtReqLoc_7 <= 6'h0;
            end
            if(_zz_366[8]) begin
              cntCmtReqLoc_8 <= 6'h0;
            end
            if(_zz_366[9]) begin
              cntCmtReqLoc_9 <= 6'h0;
            end
            if(_zz_366[10]) begin
              cntCmtReqLoc_10 <= 6'h0;
            end
            if(_zz_366[11]) begin
              cntCmtReqLoc_11 <= 6'h0;
            end
            if(_zz_366[12]) begin
              cntCmtReqLoc_12 <= 6'h0;
            end
            if(_zz_366[13]) begin
              cntCmtReqLoc_13 <= 6'h0;
            end
            if(_zz_366[14]) begin
              cntCmtReqLoc_14 <= 6'h0;
            end
            if(_zz_366[15]) begin
              cntCmtReqLoc_15 <= 6'h0;
            end
            if(_zz_366[16]) begin
              cntCmtReqLoc_16 <= 6'h0;
            end
            if(_zz_366[17]) begin
              cntCmtReqLoc_17 <= 6'h0;
            end
            if(_zz_366[18]) begin
              cntCmtReqLoc_18 <= 6'h0;
            end
            if(_zz_366[19]) begin
              cntCmtReqLoc_19 <= 6'h0;
            end
            if(_zz_366[20]) begin
              cntCmtReqLoc_20 <= 6'h0;
            end
            if(_zz_366[21]) begin
              cntCmtReqLoc_21 <= 6'h0;
            end
            if(_zz_366[22]) begin
              cntCmtReqLoc_22 <= 6'h0;
            end
            if(_zz_366[23]) begin
              cntCmtReqLoc_23 <= 6'h0;
            end
            if(_zz_366[24]) begin
              cntCmtReqLoc_24 <= 6'h0;
            end
            if(_zz_366[25]) begin
              cntCmtReqLoc_25 <= 6'h0;
            end
            if(_zz_366[26]) begin
              cntCmtReqLoc_26 <= 6'h0;
            end
            if(_zz_366[27]) begin
              cntCmtReqLoc_27 <= 6'h0;
            end
            if(_zz_366[28]) begin
              cntCmtReqLoc_28 <= 6'h0;
            end
            if(_zz_366[29]) begin
              cntCmtReqLoc_29 <= 6'h0;
            end
            if(_zz_366[30]) begin
              cntCmtReqLoc_30 <= 6'h0;
            end
            if(_zz_366[31]) begin
              cntCmtReqLoc_31 <= 6'h0;
            end
            if(_zz_366[32]) begin
              cntCmtReqLoc_32 <= 6'h0;
            end
            if(_zz_366[33]) begin
              cntCmtReqLoc_33 <= 6'h0;
            end
            if(_zz_366[34]) begin
              cntCmtReqLoc_34 <= 6'h0;
            end
            if(_zz_366[35]) begin
              cntCmtReqLoc_35 <= 6'h0;
            end
            if(_zz_366[36]) begin
              cntCmtReqLoc_36 <= 6'h0;
            end
            if(_zz_366[37]) begin
              cntCmtReqLoc_37 <= 6'h0;
            end
            if(_zz_366[38]) begin
              cntCmtReqLoc_38 <= 6'h0;
            end
            if(_zz_366[39]) begin
              cntCmtReqLoc_39 <= 6'h0;
            end
            if(_zz_366[40]) begin
              cntCmtReqLoc_40 <= 6'h0;
            end
            if(_zz_366[41]) begin
              cntCmtReqLoc_41 <= 6'h0;
            end
            if(_zz_366[42]) begin
              cntCmtReqLoc_42 <= 6'h0;
            end
            if(_zz_366[43]) begin
              cntCmtReqLoc_43 <= 6'h0;
            end
            if(_zz_366[44]) begin
              cntCmtReqLoc_44 <= 6'h0;
            end
            if(_zz_366[45]) begin
              cntCmtReqLoc_45 <= 6'h0;
            end
            if(_zz_366[46]) begin
              cntCmtReqLoc_46 <= 6'h0;
            end
            if(_zz_366[47]) begin
              cntCmtReqLoc_47 <= 6'h0;
            end
            if(_zz_366[48]) begin
              cntCmtReqLoc_48 <= 6'h0;
            end
            if(_zz_366[49]) begin
              cntCmtReqLoc_49 <= 6'h0;
            end
            if(_zz_366[50]) begin
              cntCmtReqLoc_50 <= 6'h0;
            end
            if(_zz_366[51]) begin
              cntCmtReqLoc_51 <= 6'h0;
            end
            if(_zz_366[52]) begin
              cntCmtReqLoc_52 <= 6'h0;
            end
            if(_zz_366[53]) begin
              cntCmtReqLoc_53 <= 6'h0;
            end
            if(_zz_366[54]) begin
              cntCmtReqLoc_54 <= 6'h0;
            end
            if(_zz_366[55]) begin
              cntCmtReqLoc_55 <= 6'h0;
            end
            if(_zz_366[56]) begin
              cntCmtReqLoc_56 <= 6'h0;
            end
            if(_zz_366[57]) begin
              cntCmtReqLoc_57 <= 6'h0;
            end
            if(_zz_366[58]) begin
              cntCmtReqLoc_58 <= 6'h0;
            end
            if(_zz_366[59]) begin
              cntCmtReqLoc_59 <= 6'h0;
            end
            if(_zz_366[60]) begin
              cntCmtReqLoc_60 <= 6'h0;
            end
            if(_zz_366[61]) begin
              cntCmtReqLoc_61 <= 6'h0;
            end
            if(_zz_366[62]) begin
              cntCmtReqLoc_62 <= 6'h0;
            end
            if(_zz_366[63]) begin
              cntCmtReqLoc_63 <= 6'h0;
            end
            if(_zz_367[0]) begin
              cntCmtReqRmt_0 <= 6'h0;
            end
            if(_zz_367[1]) begin
              cntCmtReqRmt_1 <= 6'h0;
            end
            if(_zz_367[2]) begin
              cntCmtReqRmt_2 <= 6'h0;
            end
            if(_zz_367[3]) begin
              cntCmtReqRmt_3 <= 6'h0;
            end
            if(_zz_367[4]) begin
              cntCmtReqRmt_4 <= 6'h0;
            end
            if(_zz_367[5]) begin
              cntCmtReqRmt_5 <= 6'h0;
            end
            if(_zz_367[6]) begin
              cntCmtReqRmt_6 <= 6'h0;
            end
            if(_zz_367[7]) begin
              cntCmtReqRmt_7 <= 6'h0;
            end
            if(_zz_367[8]) begin
              cntCmtReqRmt_8 <= 6'h0;
            end
            if(_zz_367[9]) begin
              cntCmtReqRmt_9 <= 6'h0;
            end
            if(_zz_367[10]) begin
              cntCmtReqRmt_10 <= 6'h0;
            end
            if(_zz_367[11]) begin
              cntCmtReqRmt_11 <= 6'h0;
            end
            if(_zz_367[12]) begin
              cntCmtReqRmt_12 <= 6'h0;
            end
            if(_zz_367[13]) begin
              cntCmtReqRmt_13 <= 6'h0;
            end
            if(_zz_367[14]) begin
              cntCmtReqRmt_14 <= 6'h0;
            end
            if(_zz_367[15]) begin
              cntCmtReqRmt_15 <= 6'h0;
            end
            if(_zz_367[16]) begin
              cntCmtReqRmt_16 <= 6'h0;
            end
            if(_zz_367[17]) begin
              cntCmtReqRmt_17 <= 6'h0;
            end
            if(_zz_367[18]) begin
              cntCmtReqRmt_18 <= 6'h0;
            end
            if(_zz_367[19]) begin
              cntCmtReqRmt_19 <= 6'h0;
            end
            if(_zz_367[20]) begin
              cntCmtReqRmt_20 <= 6'h0;
            end
            if(_zz_367[21]) begin
              cntCmtReqRmt_21 <= 6'h0;
            end
            if(_zz_367[22]) begin
              cntCmtReqRmt_22 <= 6'h0;
            end
            if(_zz_367[23]) begin
              cntCmtReqRmt_23 <= 6'h0;
            end
            if(_zz_367[24]) begin
              cntCmtReqRmt_24 <= 6'h0;
            end
            if(_zz_367[25]) begin
              cntCmtReqRmt_25 <= 6'h0;
            end
            if(_zz_367[26]) begin
              cntCmtReqRmt_26 <= 6'h0;
            end
            if(_zz_367[27]) begin
              cntCmtReqRmt_27 <= 6'h0;
            end
            if(_zz_367[28]) begin
              cntCmtReqRmt_28 <= 6'h0;
            end
            if(_zz_367[29]) begin
              cntCmtReqRmt_29 <= 6'h0;
            end
            if(_zz_367[30]) begin
              cntCmtReqRmt_30 <= 6'h0;
            end
            if(_zz_367[31]) begin
              cntCmtReqRmt_31 <= 6'h0;
            end
            if(_zz_367[32]) begin
              cntCmtReqRmt_32 <= 6'h0;
            end
            if(_zz_367[33]) begin
              cntCmtReqRmt_33 <= 6'h0;
            end
            if(_zz_367[34]) begin
              cntCmtReqRmt_34 <= 6'h0;
            end
            if(_zz_367[35]) begin
              cntCmtReqRmt_35 <= 6'h0;
            end
            if(_zz_367[36]) begin
              cntCmtReqRmt_36 <= 6'h0;
            end
            if(_zz_367[37]) begin
              cntCmtReqRmt_37 <= 6'h0;
            end
            if(_zz_367[38]) begin
              cntCmtReqRmt_38 <= 6'h0;
            end
            if(_zz_367[39]) begin
              cntCmtReqRmt_39 <= 6'h0;
            end
            if(_zz_367[40]) begin
              cntCmtReqRmt_40 <= 6'h0;
            end
            if(_zz_367[41]) begin
              cntCmtReqRmt_41 <= 6'h0;
            end
            if(_zz_367[42]) begin
              cntCmtReqRmt_42 <= 6'h0;
            end
            if(_zz_367[43]) begin
              cntCmtReqRmt_43 <= 6'h0;
            end
            if(_zz_367[44]) begin
              cntCmtReqRmt_44 <= 6'h0;
            end
            if(_zz_367[45]) begin
              cntCmtReqRmt_45 <= 6'h0;
            end
            if(_zz_367[46]) begin
              cntCmtReqRmt_46 <= 6'h0;
            end
            if(_zz_367[47]) begin
              cntCmtReqRmt_47 <= 6'h0;
            end
            if(_zz_367[48]) begin
              cntCmtReqRmt_48 <= 6'h0;
            end
            if(_zz_367[49]) begin
              cntCmtReqRmt_49 <= 6'h0;
            end
            if(_zz_367[50]) begin
              cntCmtReqRmt_50 <= 6'h0;
            end
            if(_zz_367[51]) begin
              cntCmtReqRmt_51 <= 6'h0;
            end
            if(_zz_367[52]) begin
              cntCmtReqRmt_52 <= 6'h0;
            end
            if(_zz_367[53]) begin
              cntCmtReqRmt_53 <= 6'h0;
            end
            if(_zz_367[54]) begin
              cntCmtReqRmt_54 <= 6'h0;
            end
            if(_zz_367[55]) begin
              cntCmtReqRmt_55 <= 6'h0;
            end
            if(_zz_367[56]) begin
              cntCmtReqRmt_56 <= 6'h0;
            end
            if(_zz_367[57]) begin
              cntCmtReqRmt_57 <= 6'h0;
            end
            if(_zz_367[58]) begin
              cntCmtReqRmt_58 <= 6'h0;
            end
            if(_zz_367[59]) begin
              cntCmtReqRmt_59 <= 6'h0;
            end
            if(_zz_367[60]) begin
              cntCmtReqRmt_60 <= 6'h0;
            end
            if(_zz_367[61]) begin
              cntCmtReqRmt_61 <= 6'h0;
            end
            if(_zz_367[62]) begin
              cntCmtReqRmt_62 <= 6'h0;
            end
            if(_zz_367[63]) begin
              cntCmtReqRmt_63 <= 6'h0;
            end
            if(_zz_368[0]) begin
              cntCmtRespLoc_0 <= 6'h0;
            end
            if(_zz_368[1]) begin
              cntCmtRespLoc_1 <= 6'h0;
            end
            if(_zz_368[2]) begin
              cntCmtRespLoc_2 <= 6'h0;
            end
            if(_zz_368[3]) begin
              cntCmtRespLoc_3 <= 6'h0;
            end
            if(_zz_368[4]) begin
              cntCmtRespLoc_4 <= 6'h0;
            end
            if(_zz_368[5]) begin
              cntCmtRespLoc_5 <= 6'h0;
            end
            if(_zz_368[6]) begin
              cntCmtRespLoc_6 <= 6'h0;
            end
            if(_zz_368[7]) begin
              cntCmtRespLoc_7 <= 6'h0;
            end
            if(_zz_368[8]) begin
              cntCmtRespLoc_8 <= 6'h0;
            end
            if(_zz_368[9]) begin
              cntCmtRespLoc_9 <= 6'h0;
            end
            if(_zz_368[10]) begin
              cntCmtRespLoc_10 <= 6'h0;
            end
            if(_zz_368[11]) begin
              cntCmtRespLoc_11 <= 6'h0;
            end
            if(_zz_368[12]) begin
              cntCmtRespLoc_12 <= 6'h0;
            end
            if(_zz_368[13]) begin
              cntCmtRespLoc_13 <= 6'h0;
            end
            if(_zz_368[14]) begin
              cntCmtRespLoc_14 <= 6'h0;
            end
            if(_zz_368[15]) begin
              cntCmtRespLoc_15 <= 6'h0;
            end
            if(_zz_368[16]) begin
              cntCmtRespLoc_16 <= 6'h0;
            end
            if(_zz_368[17]) begin
              cntCmtRespLoc_17 <= 6'h0;
            end
            if(_zz_368[18]) begin
              cntCmtRespLoc_18 <= 6'h0;
            end
            if(_zz_368[19]) begin
              cntCmtRespLoc_19 <= 6'h0;
            end
            if(_zz_368[20]) begin
              cntCmtRespLoc_20 <= 6'h0;
            end
            if(_zz_368[21]) begin
              cntCmtRespLoc_21 <= 6'h0;
            end
            if(_zz_368[22]) begin
              cntCmtRespLoc_22 <= 6'h0;
            end
            if(_zz_368[23]) begin
              cntCmtRespLoc_23 <= 6'h0;
            end
            if(_zz_368[24]) begin
              cntCmtRespLoc_24 <= 6'h0;
            end
            if(_zz_368[25]) begin
              cntCmtRespLoc_25 <= 6'h0;
            end
            if(_zz_368[26]) begin
              cntCmtRespLoc_26 <= 6'h0;
            end
            if(_zz_368[27]) begin
              cntCmtRespLoc_27 <= 6'h0;
            end
            if(_zz_368[28]) begin
              cntCmtRespLoc_28 <= 6'h0;
            end
            if(_zz_368[29]) begin
              cntCmtRespLoc_29 <= 6'h0;
            end
            if(_zz_368[30]) begin
              cntCmtRespLoc_30 <= 6'h0;
            end
            if(_zz_368[31]) begin
              cntCmtRespLoc_31 <= 6'h0;
            end
            if(_zz_368[32]) begin
              cntCmtRespLoc_32 <= 6'h0;
            end
            if(_zz_368[33]) begin
              cntCmtRespLoc_33 <= 6'h0;
            end
            if(_zz_368[34]) begin
              cntCmtRespLoc_34 <= 6'h0;
            end
            if(_zz_368[35]) begin
              cntCmtRespLoc_35 <= 6'h0;
            end
            if(_zz_368[36]) begin
              cntCmtRespLoc_36 <= 6'h0;
            end
            if(_zz_368[37]) begin
              cntCmtRespLoc_37 <= 6'h0;
            end
            if(_zz_368[38]) begin
              cntCmtRespLoc_38 <= 6'h0;
            end
            if(_zz_368[39]) begin
              cntCmtRespLoc_39 <= 6'h0;
            end
            if(_zz_368[40]) begin
              cntCmtRespLoc_40 <= 6'h0;
            end
            if(_zz_368[41]) begin
              cntCmtRespLoc_41 <= 6'h0;
            end
            if(_zz_368[42]) begin
              cntCmtRespLoc_42 <= 6'h0;
            end
            if(_zz_368[43]) begin
              cntCmtRespLoc_43 <= 6'h0;
            end
            if(_zz_368[44]) begin
              cntCmtRespLoc_44 <= 6'h0;
            end
            if(_zz_368[45]) begin
              cntCmtRespLoc_45 <= 6'h0;
            end
            if(_zz_368[46]) begin
              cntCmtRespLoc_46 <= 6'h0;
            end
            if(_zz_368[47]) begin
              cntCmtRespLoc_47 <= 6'h0;
            end
            if(_zz_368[48]) begin
              cntCmtRespLoc_48 <= 6'h0;
            end
            if(_zz_368[49]) begin
              cntCmtRespLoc_49 <= 6'h0;
            end
            if(_zz_368[50]) begin
              cntCmtRespLoc_50 <= 6'h0;
            end
            if(_zz_368[51]) begin
              cntCmtRespLoc_51 <= 6'h0;
            end
            if(_zz_368[52]) begin
              cntCmtRespLoc_52 <= 6'h0;
            end
            if(_zz_368[53]) begin
              cntCmtRespLoc_53 <= 6'h0;
            end
            if(_zz_368[54]) begin
              cntCmtRespLoc_54 <= 6'h0;
            end
            if(_zz_368[55]) begin
              cntCmtRespLoc_55 <= 6'h0;
            end
            if(_zz_368[56]) begin
              cntCmtRespLoc_56 <= 6'h0;
            end
            if(_zz_368[57]) begin
              cntCmtRespLoc_57 <= 6'h0;
            end
            if(_zz_368[58]) begin
              cntCmtRespLoc_58 <= 6'h0;
            end
            if(_zz_368[59]) begin
              cntCmtRespLoc_59 <= 6'h0;
            end
            if(_zz_368[60]) begin
              cntCmtRespLoc_60 <= 6'h0;
            end
            if(_zz_368[61]) begin
              cntCmtRespLoc_61 <= 6'h0;
            end
            if(_zz_368[62]) begin
              cntCmtRespLoc_62 <= 6'h0;
            end
            if(_zz_368[63]) begin
              cntCmtRespLoc_63 <= 6'h0;
            end
            if(_zz_369[0]) begin
              cntCmtRespRmt_0 <= 6'h0;
            end
            if(_zz_369[1]) begin
              cntCmtRespRmt_1 <= 6'h0;
            end
            if(_zz_369[2]) begin
              cntCmtRespRmt_2 <= 6'h0;
            end
            if(_zz_369[3]) begin
              cntCmtRespRmt_3 <= 6'h0;
            end
            if(_zz_369[4]) begin
              cntCmtRespRmt_4 <= 6'h0;
            end
            if(_zz_369[5]) begin
              cntCmtRespRmt_5 <= 6'h0;
            end
            if(_zz_369[6]) begin
              cntCmtRespRmt_6 <= 6'h0;
            end
            if(_zz_369[7]) begin
              cntCmtRespRmt_7 <= 6'h0;
            end
            if(_zz_369[8]) begin
              cntCmtRespRmt_8 <= 6'h0;
            end
            if(_zz_369[9]) begin
              cntCmtRespRmt_9 <= 6'h0;
            end
            if(_zz_369[10]) begin
              cntCmtRespRmt_10 <= 6'h0;
            end
            if(_zz_369[11]) begin
              cntCmtRespRmt_11 <= 6'h0;
            end
            if(_zz_369[12]) begin
              cntCmtRespRmt_12 <= 6'h0;
            end
            if(_zz_369[13]) begin
              cntCmtRespRmt_13 <= 6'h0;
            end
            if(_zz_369[14]) begin
              cntCmtRespRmt_14 <= 6'h0;
            end
            if(_zz_369[15]) begin
              cntCmtRespRmt_15 <= 6'h0;
            end
            if(_zz_369[16]) begin
              cntCmtRespRmt_16 <= 6'h0;
            end
            if(_zz_369[17]) begin
              cntCmtRespRmt_17 <= 6'h0;
            end
            if(_zz_369[18]) begin
              cntCmtRespRmt_18 <= 6'h0;
            end
            if(_zz_369[19]) begin
              cntCmtRespRmt_19 <= 6'h0;
            end
            if(_zz_369[20]) begin
              cntCmtRespRmt_20 <= 6'h0;
            end
            if(_zz_369[21]) begin
              cntCmtRespRmt_21 <= 6'h0;
            end
            if(_zz_369[22]) begin
              cntCmtRespRmt_22 <= 6'h0;
            end
            if(_zz_369[23]) begin
              cntCmtRespRmt_23 <= 6'h0;
            end
            if(_zz_369[24]) begin
              cntCmtRespRmt_24 <= 6'h0;
            end
            if(_zz_369[25]) begin
              cntCmtRespRmt_25 <= 6'h0;
            end
            if(_zz_369[26]) begin
              cntCmtRespRmt_26 <= 6'h0;
            end
            if(_zz_369[27]) begin
              cntCmtRespRmt_27 <= 6'h0;
            end
            if(_zz_369[28]) begin
              cntCmtRespRmt_28 <= 6'h0;
            end
            if(_zz_369[29]) begin
              cntCmtRespRmt_29 <= 6'h0;
            end
            if(_zz_369[30]) begin
              cntCmtRespRmt_30 <= 6'h0;
            end
            if(_zz_369[31]) begin
              cntCmtRespRmt_31 <= 6'h0;
            end
            if(_zz_369[32]) begin
              cntCmtRespRmt_32 <= 6'h0;
            end
            if(_zz_369[33]) begin
              cntCmtRespRmt_33 <= 6'h0;
            end
            if(_zz_369[34]) begin
              cntCmtRespRmt_34 <= 6'h0;
            end
            if(_zz_369[35]) begin
              cntCmtRespRmt_35 <= 6'h0;
            end
            if(_zz_369[36]) begin
              cntCmtRespRmt_36 <= 6'h0;
            end
            if(_zz_369[37]) begin
              cntCmtRespRmt_37 <= 6'h0;
            end
            if(_zz_369[38]) begin
              cntCmtRespRmt_38 <= 6'h0;
            end
            if(_zz_369[39]) begin
              cntCmtRespRmt_39 <= 6'h0;
            end
            if(_zz_369[40]) begin
              cntCmtRespRmt_40 <= 6'h0;
            end
            if(_zz_369[41]) begin
              cntCmtRespRmt_41 <= 6'h0;
            end
            if(_zz_369[42]) begin
              cntCmtRespRmt_42 <= 6'h0;
            end
            if(_zz_369[43]) begin
              cntCmtRespRmt_43 <= 6'h0;
            end
            if(_zz_369[44]) begin
              cntCmtRespRmt_44 <= 6'h0;
            end
            if(_zz_369[45]) begin
              cntCmtRespRmt_45 <= 6'h0;
            end
            if(_zz_369[46]) begin
              cntCmtRespRmt_46 <= 6'h0;
            end
            if(_zz_369[47]) begin
              cntCmtRespRmt_47 <= 6'h0;
            end
            if(_zz_369[48]) begin
              cntCmtRespRmt_48 <= 6'h0;
            end
            if(_zz_369[49]) begin
              cntCmtRespRmt_49 <= 6'h0;
            end
            if(_zz_369[50]) begin
              cntCmtRespRmt_50 <= 6'h0;
            end
            if(_zz_369[51]) begin
              cntCmtRespRmt_51 <= 6'h0;
            end
            if(_zz_369[52]) begin
              cntCmtRespRmt_52 <= 6'h0;
            end
            if(_zz_369[53]) begin
              cntCmtRespRmt_53 <= 6'h0;
            end
            if(_zz_369[54]) begin
              cntCmtRespRmt_54 <= 6'h0;
            end
            if(_zz_369[55]) begin
              cntCmtRespRmt_55 <= 6'h0;
            end
            if(_zz_369[56]) begin
              cntCmtRespRmt_56 <= 6'h0;
            end
            if(_zz_369[57]) begin
              cntCmtRespRmt_57 <= 6'h0;
            end
            if(_zz_369[58]) begin
              cntCmtRespRmt_58 <= 6'h0;
            end
            if(_zz_369[59]) begin
              cntCmtRespRmt_59 <= 6'h0;
            end
            if(_zz_369[60]) begin
              cntCmtRespRmt_60 <= 6'h0;
            end
            if(_zz_369[61]) begin
              cntCmtRespRmt_61 <= 6'h0;
            end
            if(_zz_369[62]) begin
              cntCmtRespRmt_62 <= 6'h0;
            end
            if(_zz_369[63]) begin
              cntCmtRespRmt_63 <= 6'h0;
            end
            if(_zz_370[0]) begin
              cntRlseReqLoc_0 <= 6'h0;
            end
            if(_zz_370[1]) begin
              cntRlseReqLoc_1 <= 6'h0;
            end
            if(_zz_370[2]) begin
              cntRlseReqLoc_2 <= 6'h0;
            end
            if(_zz_370[3]) begin
              cntRlseReqLoc_3 <= 6'h0;
            end
            if(_zz_370[4]) begin
              cntRlseReqLoc_4 <= 6'h0;
            end
            if(_zz_370[5]) begin
              cntRlseReqLoc_5 <= 6'h0;
            end
            if(_zz_370[6]) begin
              cntRlseReqLoc_6 <= 6'h0;
            end
            if(_zz_370[7]) begin
              cntRlseReqLoc_7 <= 6'h0;
            end
            if(_zz_370[8]) begin
              cntRlseReqLoc_8 <= 6'h0;
            end
            if(_zz_370[9]) begin
              cntRlseReqLoc_9 <= 6'h0;
            end
            if(_zz_370[10]) begin
              cntRlseReqLoc_10 <= 6'h0;
            end
            if(_zz_370[11]) begin
              cntRlseReqLoc_11 <= 6'h0;
            end
            if(_zz_370[12]) begin
              cntRlseReqLoc_12 <= 6'h0;
            end
            if(_zz_370[13]) begin
              cntRlseReqLoc_13 <= 6'h0;
            end
            if(_zz_370[14]) begin
              cntRlseReqLoc_14 <= 6'h0;
            end
            if(_zz_370[15]) begin
              cntRlseReqLoc_15 <= 6'h0;
            end
            if(_zz_370[16]) begin
              cntRlseReqLoc_16 <= 6'h0;
            end
            if(_zz_370[17]) begin
              cntRlseReqLoc_17 <= 6'h0;
            end
            if(_zz_370[18]) begin
              cntRlseReqLoc_18 <= 6'h0;
            end
            if(_zz_370[19]) begin
              cntRlseReqLoc_19 <= 6'h0;
            end
            if(_zz_370[20]) begin
              cntRlseReqLoc_20 <= 6'h0;
            end
            if(_zz_370[21]) begin
              cntRlseReqLoc_21 <= 6'h0;
            end
            if(_zz_370[22]) begin
              cntRlseReqLoc_22 <= 6'h0;
            end
            if(_zz_370[23]) begin
              cntRlseReqLoc_23 <= 6'h0;
            end
            if(_zz_370[24]) begin
              cntRlseReqLoc_24 <= 6'h0;
            end
            if(_zz_370[25]) begin
              cntRlseReqLoc_25 <= 6'h0;
            end
            if(_zz_370[26]) begin
              cntRlseReqLoc_26 <= 6'h0;
            end
            if(_zz_370[27]) begin
              cntRlseReqLoc_27 <= 6'h0;
            end
            if(_zz_370[28]) begin
              cntRlseReqLoc_28 <= 6'h0;
            end
            if(_zz_370[29]) begin
              cntRlseReqLoc_29 <= 6'h0;
            end
            if(_zz_370[30]) begin
              cntRlseReqLoc_30 <= 6'h0;
            end
            if(_zz_370[31]) begin
              cntRlseReqLoc_31 <= 6'h0;
            end
            if(_zz_370[32]) begin
              cntRlseReqLoc_32 <= 6'h0;
            end
            if(_zz_370[33]) begin
              cntRlseReqLoc_33 <= 6'h0;
            end
            if(_zz_370[34]) begin
              cntRlseReqLoc_34 <= 6'h0;
            end
            if(_zz_370[35]) begin
              cntRlseReqLoc_35 <= 6'h0;
            end
            if(_zz_370[36]) begin
              cntRlseReqLoc_36 <= 6'h0;
            end
            if(_zz_370[37]) begin
              cntRlseReqLoc_37 <= 6'h0;
            end
            if(_zz_370[38]) begin
              cntRlseReqLoc_38 <= 6'h0;
            end
            if(_zz_370[39]) begin
              cntRlseReqLoc_39 <= 6'h0;
            end
            if(_zz_370[40]) begin
              cntRlseReqLoc_40 <= 6'h0;
            end
            if(_zz_370[41]) begin
              cntRlseReqLoc_41 <= 6'h0;
            end
            if(_zz_370[42]) begin
              cntRlseReqLoc_42 <= 6'h0;
            end
            if(_zz_370[43]) begin
              cntRlseReqLoc_43 <= 6'h0;
            end
            if(_zz_370[44]) begin
              cntRlseReqLoc_44 <= 6'h0;
            end
            if(_zz_370[45]) begin
              cntRlseReqLoc_45 <= 6'h0;
            end
            if(_zz_370[46]) begin
              cntRlseReqLoc_46 <= 6'h0;
            end
            if(_zz_370[47]) begin
              cntRlseReqLoc_47 <= 6'h0;
            end
            if(_zz_370[48]) begin
              cntRlseReqLoc_48 <= 6'h0;
            end
            if(_zz_370[49]) begin
              cntRlseReqLoc_49 <= 6'h0;
            end
            if(_zz_370[50]) begin
              cntRlseReqLoc_50 <= 6'h0;
            end
            if(_zz_370[51]) begin
              cntRlseReqLoc_51 <= 6'h0;
            end
            if(_zz_370[52]) begin
              cntRlseReqLoc_52 <= 6'h0;
            end
            if(_zz_370[53]) begin
              cntRlseReqLoc_53 <= 6'h0;
            end
            if(_zz_370[54]) begin
              cntRlseReqLoc_54 <= 6'h0;
            end
            if(_zz_370[55]) begin
              cntRlseReqLoc_55 <= 6'h0;
            end
            if(_zz_370[56]) begin
              cntRlseReqLoc_56 <= 6'h0;
            end
            if(_zz_370[57]) begin
              cntRlseReqLoc_57 <= 6'h0;
            end
            if(_zz_370[58]) begin
              cntRlseReqLoc_58 <= 6'h0;
            end
            if(_zz_370[59]) begin
              cntRlseReqLoc_59 <= 6'h0;
            end
            if(_zz_370[60]) begin
              cntRlseReqLoc_60 <= 6'h0;
            end
            if(_zz_370[61]) begin
              cntRlseReqLoc_61 <= 6'h0;
            end
            if(_zz_370[62]) begin
              cntRlseReqLoc_62 <= 6'h0;
            end
            if(_zz_370[63]) begin
              cntRlseReqLoc_63 <= 6'h0;
            end
            if(_zz_371[0]) begin
              cntRlseReqRmt_0 <= 6'h0;
            end
            if(_zz_371[1]) begin
              cntRlseReqRmt_1 <= 6'h0;
            end
            if(_zz_371[2]) begin
              cntRlseReqRmt_2 <= 6'h0;
            end
            if(_zz_371[3]) begin
              cntRlseReqRmt_3 <= 6'h0;
            end
            if(_zz_371[4]) begin
              cntRlseReqRmt_4 <= 6'h0;
            end
            if(_zz_371[5]) begin
              cntRlseReqRmt_5 <= 6'h0;
            end
            if(_zz_371[6]) begin
              cntRlseReqRmt_6 <= 6'h0;
            end
            if(_zz_371[7]) begin
              cntRlseReqRmt_7 <= 6'h0;
            end
            if(_zz_371[8]) begin
              cntRlseReqRmt_8 <= 6'h0;
            end
            if(_zz_371[9]) begin
              cntRlseReqRmt_9 <= 6'h0;
            end
            if(_zz_371[10]) begin
              cntRlseReqRmt_10 <= 6'h0;
            end
            if(_zz_371[11]) begin
              cntRlseReqRmt_11 <= 6'h0;
            end
            if(_zz_371[12]) begin
              cntRlseReqRmt_12 <= 6'h0;
            end
            if(_zz_371[13]) begin
              cntRlseReqRmt_13 <= 6'h0;
            end
            if(_zz_371[14]) begin
              cntRlseReqRmt_14 <= 6'h0;
            end
            if(_zz_371[15]) begin
              cntRlseReqRmt_15 <= 6'h0;
            end
            if(_zz_371[16]) begin
              cntRlseReqRmt_16 <= 6'h0;
            end
            if(_zz_371[17]) begin
              cntRlseReqRmt_17 <= 6'h0;
            end
            if(_zz_371[18]) begin
              cntRlseReqRmt_18 <= 6'h0;
            end
            if(_zz_371[19]) begin
              cntRlseReqRmt_19 <= 6'h0;
            end
            if(_zz_371[20]) begin
              cntRlseReqRmt_20 <= 6'h0;
            end
            if(_zz_371[21]) begin
              cntRlseReqRmt_21 <= 6'h0;
            end
            if(_zz_371[22]) begin
              cntRlseReqRmt_22 <= 6'h0;
            end
            if(_zz_371[23]) begin
              cntRlseReqRmt_23 <= 6'h0;
            end
            if(_zz_371[24]) begin
              cntRlseReqRmt_24 <= 6'h0;
            end
            if(_zz_371[25]) begin
              cntRlseReqRmt_25 <= 6'h0;
            end
            if(_zz_371[26]) begin
              cntRlseReqRmt_26 <= 6'h0;
            end
            if(_zz_371[27]) begin
              cntRlseReqRmt_27 <= 6'h0;
            end
            if(_zz_371[28]) begin
              cntRlseReqRmt_28 <= 6'h0;
            end
            if(_zz_371[29]) begin
              cntRlseReqRmt_29 <= 6'h0;
            end
            if(_zz_371[30]) begin
              cntRlseReqRmt_30 <= 6'h0;
            end
            if(_zz_371[31]) begin
              cntRlseReqRmt_31 <= 6'h0;
            end
            if(_zz_371[32]) begin
              cntRlseReqRmt_32 <= 6'h0;
            end
            if(_zz_371[33]) begin
              cntRlseReqRmt_33 <= 6'h0;
            end
            if(_zz_371[34]) begin
              cntRlseReqRmt_34 <= 6'h0;
            end
            if(_zz_371[35]) begin
              cntRlseReqRmt_35 <= 6'h0;
            end
            if(_zz_371[36]) begin
              cntRlseReqRmt_36 <= 6'h0;
            end
            if(_zz_371[37]) begin
              cntRlseReqRmt_37 <= 6'h0;
            end
            if(_zz_371[38]) begin
              cntRlseReqRmt_38 <= 6'h0;
            end
            if(_zz_371[39]) begin
              cntRlseReqRmt_39 <= 6'h0;
            end
            if(_zz_371[40]) begin
              cntRlseReqRmt_40 <= 6'h0;
            end
            if(_zz_371[41]) begin
              cntRlseReqRmt_41 <= 6'h0;
            end
            if(_zz_371[42]) begin
              cntRlseReqRmt_42 <= 6'h0;
            end
            if(_zz_371[43]) begin
              cntRlseReqRmt_43 <= 6'h0;
            end
            if(_zz_371[44]) begin
              cntRlseReqRmt_44 <= 6'h0;
            end
            if(_zz_371[45]) begin
              cntRlseReqRmt_45 <= 6'h0;
            end
            if(_zz_371[46]) begin
              cntRlseReqRmt_46 <= 6'h0;
            end
            if(_zz_371[47]) begin
              cntRlseReqRmt_47 <= 6'h0;
            end
            if(_zz_371[48]) begin
              cntRlseReqRmt_48 <= 6'h0;
            end
            if(_zz_371[49]) begin
              cntRlseReqRmt_49 <= 6'h0;
            end
            if(_zz_371[50]) begin
              cntRlseReqRmt_50 <= 6'h0;
            end
            if(_zz_371[51]) begin
              cntRlseReqRmt_51 <= 6'h0;
            end
            if(_zz_371[52]) begin
              cntRlseReqRmt_52 <= 6'h0;
            end
            if(_zz_371[53]) begin
              cntRlseReqRmt_53 <= 6'h0;
            end
            if(_zz_371[54]) begin
              cntRlseReqRmt_54 <= 6'h0;
            end
            if(_zz_371[55]) begin
              cntRlseReqRmt_55 <= 6'h0;
            end
            if(_zz_371[56]) begin
              cntRlseReqRmt_56 <= 6'h0;
            end
            if(_zz_371[57]) begin
              cntRlseReqRmt_57 <= 6'h0;
            end
            if(_zz_371[58]) begin
              cntRlseReqRmt_58 <= 6'h0;
            end
            if(_zz_371[59]) begin
              cntRlseReqRmt_59 <= 6'h0;
            end
            if(_zz_371[60]) begin
              cntRlseReqRmt_60 <= 6'h0;
            end
            if(_zz_371[61]) begin
              cntRlseReqRmt_61 <= 6'h0;
            end
            if(_zz_371[62]) begin
              cntRlseReqRmt_62 <= 6'h0;
            end
            if(_zz_371[63]) begin
              cntRlseReqRmt_63 <= 6'h0;
            end
            if(_zz_372[0]) begin
              cntRlseReqWrLoc_0 <= 6'h0;
            end
            if(_zz_372[1]) begin
              cntRlseReqWrLoc_1 <= 6'h0;
            end
            if(_zz_372[2]) begin
              cntRlseReqWrLoc_2 <= 6'h0;
            end
            if(_zz_372[3]) begin
              cntRlseReqWrLoc_3 <= 6'h0;
            end
            if(_zz_372[4]) begin
              cntRlseReqWrLoc_4 <= 6'h0;
            end
            if(_zz_372[5]) begin
              cntRlseReqWrLoc_5 <= 6'h0;
            end
            if(_zz_372[6]) begin
              cntRlseReqWrLoc_6 <= 6'h0;
            end
            if(_zz_372[7]) begin
              cntRlseReqWrLoc_7 <= 6'h0;
            end
            if(_zz_372[8]) begin
              cntRlseReqWrLoc_8 <= 6'h0;
            end
            if(_zz_372[9]) begin
              cntRlseReqWrLoc_9 <= 6'h0;
            end
            if(_zz_372[10]) begin
              cntRlseReqWrLoc_10 <= 6'h0;
            end
            if(_zz_372[11]) begin
              cntRlseReqWrLoc_11 <= 6'h0;
            end
            if(_zz_372[12]) begin
              cntRlseReqWrLoc_12 <= 6'h0;
            end
            if(_zz_372[13]) begin
              cntRlseReqWrLoc_13 <= 6'h0;
            end
            if(_zz_372[14]) begin
              cntRlseReqWrLoc_14 <= 6'h0;
            end
            if(_zz_372[15]) begin
              cntRlseReqWrLoc_15 <= 6'h0;
            end
            if(_zz_372[16]) begin
              cntRlseReqWrLoc_16 <= 6'h0;
            end
            if(_zz_372[17]) begin
              cntRlseReqWrLoc_17 <= 6'h0;
            end
            if(_zz_372[18]) begin
              cntRlseReqWrLoc_18 <= 6'h0;
            end
            if(_zz_372[19]) begin
              cntRlseReqWrLoc_19 <= 6'h0;
            end
            if(_zz_372[20]) begin
              cntRlseReqWrLoc_20 <= 6'h0;
            end
            if(_zz_372[21]) begin
              cntRlseReqWrLoc_21 <= 6'h0;
            end
            if(_zz_372[22]) begin
              cntRlseReqWrLoc_22 <= 6'h0;
            end
            if(_zz_372[23]) begin
              cntRlseReqWrLoc_23 <= 6'h0;
            end
            if(_zz_372[24]) begin
              cntRlseReqWrLoc_24 <= 6'h0;
            end
            if(_zz_372[25]) begin
              cntRlseReqWrLoc_25 <= 6'h0;
            end
            if(_zz_372[26]) begin
              cntRlseReqWrLoc_26 <= 6'h0;
            end
            if(_zz_372[27]) begin
              cntRlseReqWrLoc_27 <= 6'h0;
            end
            if(_zz_372[28]) begin
              cntRlseReqWrLoc_28 <= 6'h0;
            end
            if(_zz_372[29]) begin
              cntRlseReqWrLoc_29 <= 6'h0;
            end
            if(_zz_372[30]) begin
              cntRlseReqWrLoc_30 <= 6'h0;
            end
            if(_zz_372[31]) begin
              cntRlseReqWrLoc_31 <= 6'h0;
            end
            if(_zz_372[32]) begin
              cntRlseReqWrLoc_32 <= 6'h0;
            end
            if(_zz_372[33]) begin
              cntRlseReqWrLoc_33 <= 6'h0;
            end
            if(_zz_372[34]) begin
              cntRlseReqWrLoc_34 <= 6'h0;
            end
            if(_zz_372[35]) begin
              cntRlseReqWrLoc_35 <= 6'h0;
            end
            if(_zz_372[36]) begin
              cntRlseReqWrLoc_36 <= 6'h0;
            end
            if(_zz_372[37]) begin
              cntRlseReqWrLoc_37 <= 6'h0;
            end
            if(_zz_372[38]) begin
              cntRlseReqWrLoc_38 <= 6'h0;
            end
            if(_zz_372[39]) begin
              cntRlseReqWrLoc_39 <= 6'h0;
            end
            if(_zz_372[40]) begin
              cntRlseReqWrLoc_40 <= 6'h0;
            end
            if(_zz_372[41]) begin
              cntRlseReqWrLoc_41 <= 6'h0;
            end
            if(_zz_372[42]) begin
              cntRlseReqWrLoc_42 <= 6'h0;
            end
            if(_zz_372[43]) begin
              cntRlseReqWrLoc_43 <= 6'h0;
            end
            if(_zz_372[44]) begin
              cntRlseReqWrLoc_44 <= 6'h0;
            end
            if(_zz_372[45]) begin
              cntRlseReqWrLoc_45 <= 6'h0;
            end
            if(_zz_372[46]) begin
              cntRlseReqWrLoc_46 <= 6'h0;
            end
            if(_zz_372[47]) begin
              cntRlseReqWrLoc_47 <= 6'h0;
            end
            if(_zz_372[48]) begin
              cntRlseReqWrLoc_48 <= 6'h0;
            end
            if(_zz_372[49]) begin
              cntRlseReqWrLoc_49 <= 6'h0;
            end
            if(_zz_372[50]) begin
              cntRlseReqWrLoc_50 <= 6'h0;
            end
            if(_zz_372[51]) begin
              cntRlseReqWrLoc_51 <= 6'h0;
            end
            if(_zz_372[52]) begin
              cntRlseReqWrLoc_52 <= 6'h0;
            end
            if(_zz_372[53]) begin
              cntRlseReqWrLoc_53 <= 6'h0;
            end
            if(_zz_372[54]) begin
              cntRlseReqWrLoc_54 <= 6'h0;
            end
            if(_zz_372[55]) begin
              cntRlseReqWrLoc_55 <= 6'h0;
            end
            if(_zz_372[56]) begin
              cntRlseReqWrLoc_56 <= 6'h0;
            end
            if(_zz_372[57]) begin
              cntRlseReqWrLoc_57 <= 6'h0;
            end
            if(_zz_372[58]) begin
              cntRlseReqWrLoc_58 <= 6'h0;
            end
            if(_zz_372[59]) begin
              cntRlseReqWrLoc_59 <= 6'h0;
            end
            if(_zz_372[60]) begin
              cntRlseReqWrLoc_60 <= 6'h0;
            end
            if(_zz_372[61]) begin
              cntRlseReqWrLoc_61 <= 6'h0;
            end
            if(_zz_372[62]) begin
              cntRlseReqWrLoc_62 <= 6'h0;
            end
            if(_zz_372[63]) begin
              cntRlseReqWrLoc_63 <= 6'h0;
            end
            if(_zz_373[0]) begin
              cntRlseReqWrRmt_0 <= 6'h0;
            end
            if(_zz_373[1]) begin
              cntRlseReqWrRmt_1 <= 6'h0;
            end
            if(_zz_373[2]) begin
              cntRlseReqWrRmt_2 <= 6'h0;
            end
            if(_zz_373[3]) begin
              cntRlseReqWrRmt_3 <= 6'h0;
            end
            if(_zz_373[4]) begin
              cntRlseReqWrRmt_4 <= 6'h0;
            end
            if(_zz_373[5]) begin
              cntRlseReqWrRmt_5 <= 6'h0;
            end
            if(_zz_373[6]) begin
              cntRlseReqWrRmt_6 <= 6'h0;
            end
            if(_zz_373[7]) begin
              cntRlseReqWrRmt_7 <= 6'h0;
            end
            if(_zz_373[8]) begin
              cntRlseReqWrRmt_8 <= 6'h0;
            end
            if(_zz_373[9]) begin
              cntRlseReqWrRmt_9 <= 6'h0;
            end
            if(_zz_373[10]) begin
              cntRlseReqWrRmt_10 <= 6'h0;
            end
            if(_zz_373[11]) begin
              cntRlseReqWrRmt_11 <= 6'h0;
            end
            if(_zz_373[12]) begin
              cntRlseReqWrRmt_12 <= 6'h0;
            end
            if(_zz_373[13]) begin
              cntRlseReqWrRmt_13 <= 6'h0;
            end
            if(_zz_373[14]) begin
              cntRlseReqWrRmt_14 <= 6'h0;
            end
            if(_zz_373[15]) begin
              cntRlseReqWrRmt_15 <= 6'h0;
            end
            if(_zz_373[16]) begin
              cntRlseReqWrRmt_16 <= 6'h0;
            end
            if(_zz_373[17]) begin
              cntRlseReqWrRmt_17 <= 6'h0;
            end
            if(_zz_373[18]) begin
              cntRlseReqWrRmt_18 <= 6'h0;
            end
            if(_zz_373[19]) begin
              cntRlseReqWrRmt_19 <= 6'h0;
            end
            if(_zz_373[20]) begin
              cntRlseReqWrRmt_20 <= 6'h0;
            end
            if(_zz_373[21]) begin
              cntRlseReqWrRmt_21 <= 6'h0;
            end
            if(_zz_373[22]) begin
              cntRlseReqWrRmt_22 <= 6'h0;
            end
            if(_zz_373[23]) begin
              cntRlseReqWrRmt_23 <= 6'h0;
            end
            if(_zz_373[24]) begin
              cntRlseReqWrRmt_24 <= 6'h0;
            end
            if(_zz_373[25]) begin
              cntRlseReqWrRmt_25 <= 6'h0;
            end
            if(_zz_373[26]) begin
              cntRlseReqWrRmt_26 <= 6'h0;
            end
            if(_zz_373[27]) begin
              cntRlseReqWrRmt_27 <= 6'h0;
            end
            if(_zz_373[28]) begin
              cntRlseReqWrRmt_28 <= 6'h0;
            end
            if(_zz_373[29]) begin
              cntRlseReqWrRmt_29 <= 6'h0;
            end
            if(_zz_373[30]) begin
              cntRlseReqWrRmt_30 <= 6'h0;
            end
            if(_zz_373[31]) begin
              cntRlseReqWrRmt_31 <= 6'h0;
            end
            if(_zz_373[32]) begin
              cntRlseReqWrRmt_32 <= 6'h0;
            end
            if(_zz_373[33]) begin
              cntRlseReqWrRmt_33 <= 6'h0;
            end
            if(_zz_373[34]) begin
              cntRlseReqWrRmt_34 <= 6'h0;
            end
            if(_zz_373[35]) begin
              cntRlseReqWrRmt_35 <= 6'h0;
            end
            if(_zz_373[36]) begin
              cntRlseReqWrRmt_36 <= 6'h0;
            end
            if(_zz_373[37]) begin
              cntRlseReqWrRmt_37 <= 6'h0;
            end
            if(_zz_373[38]) begin
              cntRlseReqWrRmt_38 <= 6'h0;
            end
            if(_zz_373[39]) begin
              cntRlseReqWrRmt_39 <= 6'h0;
            end
            if(_zz_373[40]) begin
              cntRlseReqWrRmt_40 <= 6'h0;
            end
            if(_zz_373[41]) begin
              cntRlseReqWrRmt_41 <= 6'h0;
            end
            if(_zz_373[42]) begin
              cntRlseReqWrRmt_42 <= 6'h0;
            end
            if(_zz_373[43]) begin
              cntRlseReqWrRmt_43 <= 6'h0;
            end
            if(_zz_373[44]) begin
              cntRlseReqWrRmt_44 <= 6'h0;
            end
            if(_zz_373[45]) begin
              cntRlseReqWrRmt_45 <= 6'h0;
            end
            if(_zz_373[46]) begin
              cntRlseReqWrRmt_46 <= 6'h0;
            end
            if(_zz_373[47]) begin
              cntRlseReqWrRmt_47 <= 6'h0;
            end
            if(_zz_373[48]) begin
              cntRlseReqWrRmt_48 <= 6'h0;
            end
            if(_zz_373[49]) begin
              cntRlseReqWrRmt_49 <= 6'h0;
            end
            if(_zz_373[50]) begin
              cntRlseReqWrRmt_50 <= 6'h0;
            end
            if(_zz_373[51]) begin
              cntRlseReqWrRmt_51 <= 6'h0;
            end
            if(_zz_373[52]) begin
              cntRlseReqWrRmt_52 <= 6'h0;
            end
            if(_zz_373[53]) begin
              cntRlseReqWrRmt_53 <= 6'h0;
            end
            if(_zz_373[54]) begin
              cntRlseReqWrRmt_54 <= 6'h0;
            end
            if(_zz_373[55]) begin
              cntRlseReqWrRmt_55 <= 6'h0;
            end
            if(_zz_373[56]) begin
              cntRlseReqWrRmt_56 <= 6'h0;
            end
            if(_zz_373[57]) begin
              cntRlseReqWrRmt_57 <= 6'h0;
            end
            if(_zz_373[58]) begin
              cntRlseReqWrRmt_58 <= 6'h0;
            end
            if(_zz_373[59]) begin
              cntRlseReqWrRmt_59 <= 6'h0;
            end
            if(_zz_373[60]) begin
              cntRlseReqWrRmt_60 <= 6'h0;
            end
            if(_zz_373[61]) begin
              cntRlseReqWrRmt_61 <= 6'h0;
            end
            if(_zz_373[62]) begin
              cntRlseReqWrRmt_62 <= 6'h0;
            end
            if(_zz_373[63]) begin
              cntRlseReqWrRmt_63 <= 6'h0;
            end
            if(_zz_374[0]) begin
              cntRlseRespLoc_0 <= 6'h0;
            end
            if(_zz_374[1]) begin
              cntRlseRespLoc_1 <= 6'h0;
            end
            if(_zz_374[2]) begin
              cntRlseRespLoc_2 <= 6'h0;
            end
            if(_zz_374[3]) begin
              cntRlseRespLoc_3 <= 6'h0;
            end
            if(_zz_374[4]) begin
              cntRlseRespLoc_4 <= 6'h0;
            end
            if(_zz_374[5]) begin
              cntRlseRespLoc_5 <= 6'h0;
            end
            if(_zz_374[6]) begin
              cntRlseRespLoc_6 <= 6'h0;
            end
            if(_zz_374[7]) begin
              cntRlseRespLoc_7 <= 6'h0;
            end
            if(_zz_374[8]) begin
              cntRlseRespLoc_8 <= 6'h0;
            end
            if(_zz_374[9]) begin
              cntRlseRespLoc_9 <= 6'h0;
            end
            if(_zz_374[10]) begin
              cntRlseRespLoc_10 <= 6'h0;
            end
            if(_zz_374[11]) begin
              cntRlseRespLoc_11 <= 6'h0;
            end
            if(_zz_374[12]) begin
              cntRlseRespLoc_12 <= 6'h0;
            end
            if(_zz_374[13]) begin
              cntRlseRespLoc_13 <= 6'h0;
            end
            if(_zz_374[14]) begin
              cntRlseRespLoc_14 <= 6'h0;
            end
            if(_zz_374[15]) begin
              cntRlseRespLoc_15 <= 6'h0;
            end
            if(_zz_374[16]) begin
              cntRlseRespLoc_16 <= 6'h0;
            end
            if(_zz_374[17]) begin
              cntRlseRespLoc_17 <= 6'h0;
            end
            if(_zz_374[18]) begin
              cntRlseRespLoc_18 <= 6'h0;
            end
            if(_zz_374[19]) begin
              cntRlseRespLoc_19 <= 6'h0;
            end
            if(_zz_374[20]) begin
              cntRlseRespLoc_20 <= 6'h0;
            end
            if(_zz_374[21]) begin
              cntRlseRespLoc_21 <= 6'h0;
            end
            if(_zz_374[22]) begin
              cntRlseRespLoc_22 <= 6'h0;
            end
            if(_zz_374[23]) begin
              cntRlseRespLoc_23 <= 6'h0;
            end
            if(_zz_374[24]) begin
              cntRlseRespLoc_24 <= 6'h0;
            end
            if(_zz_374[25]) begin
              cntRlseRespLoc_25 <= 6'h0;
            end
            if(_zz_374[26]) begin
              cntRlseRespLoc_26 <= 6'h0;
            end
            if(_zz_374[27]) begin
              cntRlseRespLoc_27 <= 6'h0;
            end
            if(_zz_374[28]) begin
              cntRlseRespLoc_28 <= 6'h0;
            end
            if(_zz_374[29]) begin
              cntRlseRespLoc_29 <= 6'h0;
            end
            if(_zz_374[30]) begin
              cntRlseRespLoc_30 <= 6'h0;
            end
            if(_zz_374[31]) begin
              cntRlseRespLoc_31 <= 6'h0;
            end
            if(_zz_374[32]) begin
              cntRlseRespLoc_32 <= 6'h0;
            end
            if(_zz_374[33]) begin
              cntRlseRespLoc_33 <= 6'h0;
            end
            if(_zz_374[34]) begin
              cntRlseRespLoc_34 <= 6'h0;
            end
            if(_zz_374[35]) begin
              cntRlseRespLoc_35 <= 6'h0;
            end
            if(_zz_374[36]) begin
              cntRlseRespLoc_36 <= 6'h0;
            end
            if(_zz_374[37]) begin
              cntRlseRespLoc_37 <= 6'h0;
            end
            if(_zz_374[38]) begin
              cntRlseRespLoc_38 <= 6'h0;
            end
            if(_zz_374[39]) begin
              cntRlseRespLoc_39 <= 6'h0;
            end
            if(_zz_374[40]) begin
              cntRlseRespLoc_40 <= 6'h0;
            end
            if(_zz_374[41]) begin
              cntRlseRespLoc_41 <= 6'h0;
            end
            if(_zz_374[42]) begin
              cntRlseRespLoc_42 <= 6'h0;
            end
            if(_zz_374[43]) begin
              cntRlseRespLoc_43 <= 6'h0;
            end
            if(_zz_374[44]) begin
              cntRlseRespLoc_44 <= 6'h0;
            end
            if(_zz_374[45]) begin
              cntRlseRespLoc_45 <= 6'h0;
            end
            if(_zz_374[46]) begin
              cntRlseRespLoc_46 <= 6'h0;
            end
            if(_zz_374[47]) begin
              cntRlseRespLoc_47 <= 6'h0;
            end
            if(_zz_374[48]) begin
              cntRlseRespLoc_48 <= 6'h0;
            end
            if(_zz_374[49]) begin
              cntRlseRespLoc_49 <= 6'h0;
            end
            if(_zz_374[50]) begin
              cntRlseRespLoc_50 <= 6'h0;
            end
            if(_zz_374[51]) begin
              cntRlseRespLoc_51 <= 6'h0;
            end
            if(_zz_374[52]) begin
              cntRlseRespLoc_52 <= 6'h0;
            end
            if(_zz_374[53]) begin
              cntRlseRespLoc_53 <= 6'h0;
            end
            if(_zz_374[54]) begin
              cntRlseRespLoc_54 <= 6'h0;
            end
            if(_zz_374[55]) begin
              cntRlseRespLoc_55 <= 6'h0;
            end
            if(_zz_374[56]) begin
              cntRlseRespLoc_56 <= 6'h0;
            end
            if(_zz_374[57]) begin
              cntRlseRespLoc_57 <= 6'h0;
            end
            if(_zz_374[58]) begin
              cntRlseRespLoc_58 <= 6'h0;
            end
            if(_zz_374[59]) begin
              cntRlseRespLoc_59 <= 6'h0;
            end
            if(_zz_374[60]) begin
              cntRlseRespLoc_60 <= 6'h0;
            end
            if(_zz_374[61]) begin
              cntRlseRespLoc_61 <= 6'h0;
            end
            if(_zz_374[62]) begin
              cntRlseRespLoc_62 <= 6'h0;
            end
            if(_zz_374[63]) begin
              cntRlseRespLoc_63 <= 6'h0;
            end
            if(_zz_375[0]) begin
              cntRlseRespRmt_0 <= 6'h0;
            end
            if(_zz_375[1]) begin
              cntRlseRespRmt_1 <= 6'h0;
            end
            if(_zz_375[2]) begin
              cntRlseRespRmt_2 <= 6'h0;
            end
            if(_zz_375[3]) begin
              cntRlseRespRmt_3 <= 6'h0;
            end
            if(_zz_375[4]) begin
              cntRlseRespRmt_4 <= 6'h0;
            end
            if(_zz_375[5]) begin
              cntRlseRespRmt_5 <= 6'h0;
            end
            if(_zz_375[6]) begin
              cntRlseRespRmt_6 <= 6'h0;
            end
            if(_zz_375[7]) begin
              cntRlseRespRmt_7 <= 6'h0;
            end
            if(_zz_375[8]) begin
              cntRlseRespRmt_8 <= 6'h0;
            end
            if(_zz_375[9]) begin
              cntRlseRespRmt_9 <= 6'h0;
            end
            if(_zz_375[10]) begin
              cntRlseRespRmt_10 <= 6'h0;
            end
            if(_zz_375[11]) begin
              cntRlseRespRmt_11 <= 6'h0;
            end
            if(_zz_375[12]) begin
              cntRlseRespRmt_12 <= 6'h0;
            end
            if(_zz_375[13]) begin
              cntRlseRespRmt_13 <= 6'h0;
            end
            if(_zz_375[14]) begin
              cntRlseRespRmt_14 <= 6'h0;
            end
            if(_zz_375[15]) begin
              cntRlseRespRmt_15 <= 6'h0;
            end
            if(_zz_375[16]) begin
              cntRlseRespRmt_16 <= 6'h0;
            end
            if(_zz_375[17]) begin
              cntRlseRespRmt_17 <= 6'h0;
            end
            if(_zz_375[18]) begin
              cntRlseRespRmt_18 <= 6'h0;
            end
            if(_zz_375[19]) begin
              cntRlseRespRmt_19 <= 6'h0;
            end
            if(_zz_375[20]) begin
              cntRlseRespRmt_20 <= 6'h0;
            end
            if(_zz_375[21]) begin
              cntRlseRespRmt_21 <= 6'h0;
            end
            if(_zz_375[22]) begin
              cntRlseRespRmt_22 <= 6'h0;
            end
            if(_zz_375[23]) begin
              cntRlseRespRmt_23 <= 6'h0;
            end
            if(_zz_375[24]) begin
              cntRlseRespRmt_24 <= 6'h0;
            end
            if(_zz_375[25]) begin
              cntRlseRespRmt_25 <= 6'h0;
            end
            if(_zz_375[26]) begin
              cntRlseRespRmt_26 <= 6'h0;
            end
            if(_zz_375[27]) begin
              cntRlseRespRmt_27 <= 6'h0;
            end
            if(_zz_375[28]) begin
              cntRlseRespRmt_28 <= 6'h0;
            end
            if(_zz_375[29]) begin
              cntRlseRespRmt_29 <= 6'h0;
            end
            if(_zz_375[30]) begin
              cntRlseRespRmt_30 <= 6'h0;
            end
            if(_zz_375[31]) begin
              cntRlseRespRmt_31 <= 6'h0;
            end
            if(_zz_375[32]) begin
              cntRlseRespRmt_32 <= 6'h0;
            end
            if(_zz_375[33]) begin
              cntRlseRespRmt_33 <= 6'h0;
            end
            if(_zz_375[34]) begin
              cntRlseRespRmt_34 <= 6'h0;
            end
            if(_zz_375[35]) begin
              cntRlseRespRmt_35 <= 6'h0;
            end
            if(_zz_375[36]) begin
              cntRlseRespRmt_36 <= 6'h0;
            end
            if(_zz_375[37]) begin
              cntRlseRespRmt_37 <= 6'h0;
            end
            if(_zz_375[38]) begin
              cntRlseRespRmt_38 <= 6'h0;
            end
            if(_zz_375[39]) begin
              cntRlseRespRmt_39 <= 6'h0;
            end
            if(_zz_375[40]) begin
              cntRlseRespRmt_40 <= 6'h0;
            end
            if(_zz_375[41]) begin
              cntRlseRespRmt_41 <= 6'h0;
            end
            if(_zz_375[42]) begin
              cntRlseRespRmt_42 <= 6'h0;
            end
            if(_zz_375[43]) begin
              cntRlseRespRmt_43 <= 6'h0;
            end
            if(_zz_375[44]) begin
              cntRlseRespRmt_44 <= 6'h0;
            end
            if(_zz_375[45]) begin
              cntRlseRespRmt_45 <= 6'h0;
            end
            if(_zz_375[46]) begin
              cntRlseRespRmt_46 <= 6'h0;
            end
            if(_zz_375[47]) begin
              cntRlseRespRmt_47 <= 6'h0;
            end
            if(_zz_375[48]) begin
              cntRlseRespRmt_48 <= 6'h0;
            end
            if(_zz_375[49]) begin
              cntRlseRespRmt_49 <= 6'h0;
            end
            if(_zz_375[50]) begin
              cntRlseRespRmt_50 <= 6'h0;
            end
            if(_zz_375[51]) begin
              cntRlseRespRmt_51 <= 6'h0;
            end
            if(_zz_375[52]) begin
              cntRlseRespRmt_52 <= 6'h0;
            end
            if(_zz_375[53]) begin
              cntRlseRespRmt_53 <= 6'h0;
            end
            if(_zz_375[54]) begin
              cntRlseRespRmt_54 <= 6'h0;
            end
            if(_zz_375[55]) begin
              cntRlseRespRmt_55 <= 6'h0;
            end
            if(_zz_375[56]) begin
              cntRlseRespRmt_56 <= 6'h0;
            end
            if(_zz_375[57]) begin
              cntRlseRespRmt_57 <= 6'h0;
            end
            if(_zz_375[58]) begin
              cntRlseRespRmt_58 <= 6'h0;
            end
            if(_zz_375[59]) begin
              cntRlseRespRmt_59 <= 6'h0;
            end
            if(_zz_375[60]) begin
              cntRlseRespRmt_60 <= 6'h0;
            end
            if(_zz_375[61]) begin
              cntRlseRespRmt_61 <= 6'h0;
            end
            if(_zz_375[62]) begin
              cntRlseRespRmt_62 <= 6'h0;
            end
            if(_zz_375[63]) begin
              cntRlseRespRmt_63 <= 6'h0;
            end
            if(_zz_376[0]) begin
              cntTimeOut_0 <= 24'h0;
            end
            if(_zz_376[1]) begin
              cntTimeOut_1 <= 24'h0;
            end
            if(_zz_376[2]) begin
              cntTimeOut_2 <= 24'h0;
            end
            if(_zz_376[3]) begin
              cntTimeOut_3 <= 24'h0;
            end
            if(_zz_376[4]) begin
              cntTimeOut_4 <= 24'h0;
            end
            if(_zz_376[5]) begin
              cntTimeOut_5 <= 24'h0;
            end
            if(_zz_376[6]) begin
              cntTimeOut_6 <= 24'h0;
            end
            if(_zz_376[7]) begin
              cntTimeOut_7 <= 24'h0;
            end
            if(_zz_376[8]) begin
              cntTimeOut_8 <= 24'h0;
            end
            if(_zz_376[9]) begin
              cntTimeOut_9 <= 24'h0;
            end
            if(_zz_376[10]) begin
              cntTimeOut_10 <= 24'h0;
            end
            if(_zz_376[11]) begin
              cntTimeOut_11 <= 24'h0;
            end
            if(_zz_376[12]) begin
              cntTimeOut_12 <= 24'h0;
            end
            if(_zz_376[13]) begin
              cntTimeOut_13 <= 24'h0;
            end
            if(_zz_376[14]) begin
              cntTimeOut_14 <= 24'h0;
            end
            if(_zz_376[15]) begin
              cntTimeOut_15 <= 24'h0;
            end
            if(_zz_376[16]) begin
              cntTimeOut_16 <= 24'h0;
            end
            if(_zz_376[17]) begin
              cntTimeOut_17 <= 24'h0;
            end
            if(_zz_376[18]) begin
              cntTimeOut_18 <= 24'h0;
            end
            if(_zz_376[19]) begin
              cntTimeOut_19 <= 24'h0;
            end
            if(_zz_376[20]) begin
              cntTimeOut_20 <= 24'h0;
            end
            if(_zz_376[21]) begin
              cntTimeOut_21 <= 24'h0;
            end
            if(_zz_376[22]) begin
              cntTimeOut_22 <= 24'h0;
            end
            if(_zz_376[23]) begin
              cntTimeOut_23 <= 24'h0;
            end
            if(_zz_376[24]) begin
              cntTimeOut_24 <= 24'h0;
            end
            if(_zz_376[25]) begin
              cntTimeOut_25 <= 24'h0;
            end
            if(_zz_376[26]) begin
              cntTimeOut_26 <= 24'h0;
            end
            if(_zz_376[27]) begin
              cntTimeOut_27 <= 24'h0;
            end
            if(_zz_376[28]) begin
              cntTimeOut_28 <= 24'h0;
            end
            if(_zz_376[29]) begin
              cntTimeOut_29 <= 24'h0;
            end
            if(_zz_376[30]) begin
              cntTimeOut_30 <= 24'h0;
            end
            if(_zz_376[31]) begin
              cntTimeOut_31 <= 24'h0;
            end
            if(_zz_376[32]) begin
              cntTimeOut_32 <= 24'h0;
            end
            if(_zz_376[33]) begin
              cntTimeOut_33 <= 24'h0;
            end
            if(_zz_376[34]) begin
              cntTimeOut_34 <= 24'h0;
            end
            if(_zz_376[35]) begin
              cntTimeOut_35 <= 24'h0;
            end
            if(_zz_376[36]) begin
              cntTimeOut_36 <= 24'h0;
            end
            if(_zz_376[37]) begin
              cntTimeOut_37 <= 24'h0;
            end
            if(_zz_376[38]) begin
              cntTimeOut_38 <= 24'h0;
            end
            if(_zz_376[39]) begin
              cntTimeOut_39 <= 24'h0;
            end
            if(_zz_376[40]) begin
              cntTimeOut_40 <= 24'h0;
            end
            if(_zz_376[41]) begin
              cntTimeOut_41 <= 24'h0;
            end
            if(_zz_376[42]) begin
              cntTimeOut_42 <= 24'h0;
            end
            if(_zz_376[43]) begin
              cntTimeOut_43 <= 24'h0;
            end
            if(_zz_376[44]) begin
              cntTimeOut_44 <= 24'h0;
            end
            if(_zz_376[45]) begin
              cntTimeOut_45 <= 24'h0;
            end
            if(_zz_376[46]) begin
              cntTimeOut_46 <= 24'h0;
            end
            if(_zz_376[47]) begin
              cntTimeOut_47 <= 24'h0;
            end
            if(_zz_376[48]) begin
              cntTimeOut_48 <= 24'h0;
            end
            if(_zz_376[49]) begin
              cntTimeOut_49 <= 24'h0;
            end
            if(_zz_376[50]) begin
              cntTimeOut_50 <= 24'h0;
            end
            if(_zz_376[51]) begin
              cntTimeOut_51 <= 24'h0;
            end
            if(_zz_376[52]) begin
              cntTimeOut_52 <= 24'h0;
            end
            if(_zz_376[53]) begin
              cntTimeOut_53 <= 24'h0;
            end
            if(_zz_376[54]) begin
              cntTimeOut_54 <= 24'h0;
            end
            if(_zz_376[55]) begin
              cntTimeOut_55 <= 24'h0;
            end
            if(_zz_376[56]) begin
              cntTimeOut_56 <= 24'h0;
            end
            if(_zz_376[57]) begin
              cntTimeOut_57 <= 24'h0;
            end
            if(_zz_376[58]) begin
              cntTimeOut_58 <= 24'h0;
            end
            if(_zz_376[59]) begin
              cntTimeOut_59 <= 24'h0;
            end
            if(_zz_376[60]) begin
              cntTimeOut_60 <= 24'h0;
            end
            if(_zz_376[61]) begin
              cntTimeOut_61 <= 24'h0;
            end
            if(_zz_376[62]) begin
              cntTimeOut_62 <= 24'h0;
            end
            if(_zz_376[63]) begin
              cntTimeOut_63 <= 24'h0;
            end
            if(_zz_377[0]) begin
              rReqDone_0 <= 1'b0;
            end
            if(_zz_377[1]) begin
              rReqDone_1 <= 1'b0;
            end
            if(_zz_377[2]) begin
              rReqDone_2 <= 1'b0;
            end
            if(_zz_377[3]) begin
              rReqDone_3 <= 1'b0;
            end
            if(_zz_377[4]) begin
              rReqDone_4 <= 1'b0;
            end
            if(_zz_377[5]) begin
              rReqDone_5 <= 1'b0;
            end
            if(_zz_377[6]) begin
              rReqDone_6 <= 1'b0;
            end
            if(_zz_377[7]) begin
              rReqDone_7 <= 1'b0;
            end
            if(_zz_377[8]) begin
              rReqDone_8 <= 1'b0;
            end
            if(_zz_377[9]) begin
              rReqDone_9 <= 1'b0;
            end
            if(_zz_377[10]) begin
              rReqDone_10 <= 1'b0;
            end
            if(_zz_377[11]) begin
              rReqDone_11 <= 1'b0;
            end
            if(_zz_377[12]) begin
              rReqDone_12 <= 1'b0;
            end
            if(_zz_377[13]) begin
              rReqDone_13 <= 1'b0;
            end
            if(_zz_377[14]) begin
              rReqDone_14 <= 1'b0;
            end
            if(_zz_377[15]) begin
              rReqDone_15 <= 1'b0;
            end
            if(_zz_377[16]) begin
              rReqDone_16 <= 1'b0;
            end
            if(_zz_377[17]) begin
              rReqDone_17 <= 1'b0;
            end
            if(_zz_377[18]) begin
              rReqDone_18 <= 1'b0;
            end
            if(_zz_377[19]) begin
              rReqDone_19 <= 1'b0;
            end
            if(_zz_377[20]) begin
              rReqDone_20 <= 1'b0;
            end
            if(_zz_377[21]) begin
              rReqDone_21 <= 1'b0;
            end
            if(_zz_377[22]) begin
              rReqDone_22 <= 1'b0;
            end
            if(_zz_377[23]) begin
              rReqDone_23 <= 1'b0;
            end
            if(_zz_377[24]) begin
              rReqDone_24 <= 1'b0;
            end
            if(_zz_377[25]) begin
              rReqDone_25 <= 1'b0;
            end
            if(_zz_377[26]) begin
              rReqDone_26 <= 1'b0;
            end
            if(_zz_377[27]) begin
              rReqDone_27 <= 1'b0;
            end
            if(_zz_377[28]) begin
              rReqDone_28 <= 1'b0;
            end
            if(_zz_377[29]) begin
              rReqDone_29 <= 1'b0;
            end
            if(_zz_377[30]) begin
              rReqDone_30 <= 1'b0;
            end
            if(_zz_377[31]) begin
              rReqDone_31 <= 1'b0;
            end
            if(_zz_377[32]) begin
              rReqDone_32 <= 1'b0;
            end
            if(_zz_377[33]) begin
              rReqDone_33 <= 1'b0;
            end
            if(_zz_377[34]) begin
              rReqDone_34 <= 1'b0;
            end
            if(_zz_377[35]) begin
              rReqDone_35 <= 1'b0;
            end
            if(_zz_377[36]) begin
              rReqDone_36 <= 1'b0;
            end
            if(_zz_377[37]) begin
              rReqDone_37 <= 1'b0;
            end
            if(_zz_377[38]) begin
              rReqDone_38 <= 1'b0;
            end
            if(_zz_377[39]) begin
              rReqDone_39 <= 1'b0;
            end
            if(_zz_377[40]) begin
              rReqDone_40 <= 1'b0;
            end
            if(_zz_377[41]) begin
              rReqDone_41 <= 1'b0;
            end
            if(_zz_377[42]) begin
              rReqDone_42 <= 1'b0;
            end
            if(_zz_377[43]) begin
              rReqDone_43 <= 1'b0;
            end
            if(_zz_377[44]) begin
              rReqDone_44 <= 1'b0;
            end
            if(_zz_377[45]) begin
              rReqDone_45 <= 1'b0;
            end
            if(_zz_377[46]) begin
              rReqDone_46 <= 1'b0;
            end
            if(_zz_377[47]) begin
              rReqDone_47 <= 1'b0;
            end
            if(_zz_377[48]) begin
              rReqDone_48 <= 1'b0;
            end
            if(_zz_377[49]) begin
              rReqDone_49 <= 1'b0;
            end
            if(_zz_377[50]) begin
              rReqDone_50 <= 1'b0;
            end
            if(_zz_377[51]) begin
              rReqDone_51 <= 1'b0;
            end
            if(_zz_377[52]) begin
              rReqDone_52 <= 1'b0;
            end
            if(_zz_377[53]) begin
              rReqDone_53 <= 1'b0;
            end
            if(_zz_377[54]) begin
              rReqDone_54 <= 1'b0;
            end
            if(_zz_377[55]) begin
              rReqDone_55 <= 1'b0;
            end
            if(_zz_377[56]) begin
              rReqDone_56 <= 1'b0;
            end
            if(_zz_377[57]) begin
              rReqDone_57 <= 1'b0;
            end
            if(_zz_377[58]) begin
              rReqDone_58 <= 1'b0;
            end
            if(_zz_377[59]) begin
              rReqDone_59 <= 1'b0;
            end
            if(_zz_377[60]) begin
              rReqDone_60 <= 1'b0;
            end
            if(_zz_377[61]) begin
              rReqDone_61 <= 1'b0;
            end
            if(_zz_377[62]) begin
              rReqDone_62 <= 1'b0;
            end
            if(_zz_377[63]) begin
              rReqDone_63 <= 1'b0;
            end
            if(_zz_378[0]) begin
              rAbort_0 <= 1'b0;
            end
            if(_zz_378[1]) begin
              rAbort_1 <= 1'b0;
            end
            if(_zz_378[2]) begin
              rAbort_2 <= 1'b0;
            end
            if(_zz_378[3]) begin
              rAbort_3 <= 1'b0;
            end
            if(_zz_378[4]) begin
              rAbort_4 <= 1'b0;
            end
            if(_zz_378[5]) begin
              rAbort_5 <= 1'b0;
            end
            if(_zz_378[6]) begin
              rAbort_6 <= 1'b0;
            end
            if(_zz_378[7]) begin
              rAbort_7 <= 1'b0;
            end
            if(_zz_378[8]) begin
              rAbort_8 <= 1'b0;
            end
            if(_zz_378[9]) begin
              rAbort_9 <= 1'b0;
            end
            if(_zz_378[10]) begin
              rAbort_10 <= 1'b0;
            end
            if(_zz_378[11]) begin
              rAbort_11 <= 1'b0;
            end
            if(_zz_378[12]) begin
              rAbort_12 <= 1'b0;
            end
            if(_zz_378[13]) begin
              rAbort_13 <= 1'b0;
            end
            if(_zz_378[14]) begin
              rAbort_14 <= 1'b0;
            end
            if(_zz_378[15]) begin
              rAbort_15 <= 1'b0;
            end
            if(_zz_378[16]) begin
              rAbort_16 <= 1'b0;
            end
            if(_zz_378[17]) begin
              rAbort_17 <= 1'b0;
            end
            if(_zz_378[18]) begin
              rAbort_18 <= 1'b0;
            end
            if(_zz_378[19]) begin
              rAbort_19 <= 1'b0;
            end
            if(_zz_378[20]) begin
              rAbort_20 <= 1'b0;
            end
            if(_zz_378[21]) begin
              rAbort_21 <= 1'b0;
            end
            if(_zz_378[22]) begin
              rAbort_22 <= 1'b0;
            end
            if(_zz_378[23]) begin
              rAbort_23 <= 1'b0;
            end
            if(_zz_378[24]) begin
              rAbort_24 <= 1'b0;
            end
            if(_zz_378[25]) begin
              rAbort_25 <= 1'b0;
            end
            if(_zz_378[26]) begin
              rAbort_26 <= 1'b0;
            end
            if(_zz_378[27]) begin
              rAbort_27 <= 1'b0;
            end
            if(_zz_378[28]) begin
              rAbort_28 <= 1'b0;
            end
            if(_zz_378[29]) begin
              rAbort_29 <= 1'b0;
            end
            if(_zz_378[30]) begin
              rAbort_30 <= 1'b0;
            end
            if(_zz_378[31]) begin
              rAbort_31 <= 1'b0;
            end
            if(_zz_378[32]) begin
              rAbort_32 <= 1'b0;
            end
            if(_zz_378[33]) begin
              rAbort_33 <= 1'b0;
            end
            if(_zz_378[34]) begin
              rAbort_34 <= 1'b0;
            end
            if(_zz_378[35]) begin
              rAbort_35 <= 1'b0;
            end
            if(_zz_378[36]) begin
              rAbort_36 <= 1'b0;
            end
            if(_zz_378[37]) begin
              rAbort_37 <= 1'b0;
            end
            if(_zz_378[38]) begin
              rAbort_38 <= 1'b0;
            end
            if(_zz_378[39]) begin
              rAbort_39 <= 1'b0;
            end
            if(_zz_378[40]) begin
              rAbort_40 <= 1'b0;
            end
            if(_zz_378[41]) begin
              rAbort_41 <= 1'b0;
            end
            if(_zz_378[42]) begin
              rAbort_42 <= 1'b0;
            end
            if(_zz_378[43]) begin
              rAbort_43 <= 1'b0;
            end
            if(_zz_378[44]) begin
              rAbort_44 <= 1'b0;
            end
            if(_zz_378[45]) begin
              rAbort_45 <= 1'b0;
            end
            if(_zz_378[46]) begin
              rAbort_46 <= 1'b0;
            end
            if(_zz_378[47]) begin
              rAbort_47 <= 1'b0;
            end
            if(_zz_378[48]) begin
              rAbort_48 <= 1'b0;
            end
            if(_zz_378[49]) begin
              rAbort_49 <= 1'b0;
            end
            if(_zz_378[50]) begin
              rAbort_50 <= 1'b0;
            end
            if(_zz_378[51]) begin
              rAbort_51 <= 1'b0;
            end
            if(_zz_378[52]) begin
              rAbort_52 <= 1'b0;
            end
            if(_zz_378[53]) begin
              rAbort_53 <= 1'b0;
            end
            if(_zz_378[54]) begin
              rAbort_54 <= 1'b0;
            end
            if(_zz_378[55]) begin
              rAbort_55 <= 1'b0;
            end
            if(_zz_378[56]) begin
              rAbort_56 <= 1'b0;
            end
            if(_zz_378[57]) begin
              rAbort_57 <= 1'b0;
            end
            if(_zz_378[58]) begin
              rAbort_58 <= 1'b0;
            end
            if(_zz_378[59]) begin
              rAbort_59 <= 1'b0;
            end
            if(_zz_378[60]) begin
              rAbort_60 <= 1'b0;
            end
            if(_zz_378[61]) begin
              rAbort_61 <= 1'b0;
            end
            if(_zz_378[62]) begin
              rAbort_62 <= 1'b0;
            end
            if(_zz_378[63]) begin
              rAbort_63 <= 1'b0;
            end
            if(_zz_351[0]) begin
              rRlseDone_0 <= 1'b0;
            end
            if(_zz_351[1]) begin
              rRlseDone_1 <= 1'b0;
            end
            if(_zz_351[2]) begin
              rRlseDone_2 <= 1'b0;
            end
            if(_zz_351[3]) begin
              rRlseDone_3 <= 1'b0;
            end
            if(_zz_351[4]) begin
              rRlseDone_4 <= 1'b0;
            end
            if(_zz_351[5]) begin
              rRlseDone_5 <= 1'b0;
            end
            if(_zz_351[6]) begin
              rRlseDone_6 <= 1'b0;
            end
            if(_zz_351[7]) begin
              rRlseDone_7 <= 1'b0;
            end
            if(_zz_351[8]) begin
              rRlseDone_8 <= 1'b0;
            end
            if(_zz_351[9]) begin
              rRlseDone_9 <= 1'b0;
            end
            if(_zz_351[10]) begin
              rRlseDone_10 <= 1'b0;
            end
            if(_zz_351[11]) begin
              rRlseDone_11 <= 1'b0;
            end
            if(_zz_351[12]) begin
              rRlseDone_12 <= 1'b0;
            end
            if(_zz_351[13]) begin
              rRlseDone_13 <= 1'b0;
            end
            if(_zz_351[14]) begin
              rRlseDone_14 <= 1'b0;
            end
            if(_zz_351[15]) begin
              rRlseDone_15 <= 1'b0;
            end
            if(_zz_351[16]) begin
              rRlseDone_16 <= 1'b0;
            end
            if(_zz_351[17]) begin
              rRlseDone_17 <= 1'b0;
            end
            if(_zz_351[18]) begin
              rRlseDone_18 <= 1'b0;
            end
            if(_zz_351[19]) begin
              rRlseDone_19 <= 1'b0;
            end
            if(_zz_351[20]) begin
              rRlseDone_20 <= 1'b0;
            end
            if(_zz_351[21]) begin
              rRlseDone_21 <= 1'b0;
            end
            if(_zz_351[22]) begin
              rRlseDone_22 <= 1'b0;
            end
            if(_zz_351[23]) begin
              rRlseDone_23 <= 1'b0;
            end
            if(_zz_351[24]) begin
              rRlseDone_24 <= 1'b0;
            end
            if(_zz_351[25]) begin
              rRlseDone_25 <= 1'b0;
            end
            if(_zz_351[26]) begin
              rRlseDone_26 <= 1'b0;
            end
            if(_zz_351[27]) begin
              rRlseDone_27 <= 1'b0;
            end
            if(_zz_351[28]) begin
              rRlseDone_28 <= 1'b0;
            end
            if(_zz_351[29]) begin
              rRlseDone_29 <= 1'b0;
            end
            if(_zz_351[30]) begin
              rRlseDone_30 <= 1'b0;
            end
            if(_zz_351[31]) begin
              rRlseDone_31 <= 1'b0;
            end
            if(_zz_351[32]) begin
              rRlseDone_32 <= 1'b0;
            end
            if(_zz_351[33]) begin
              rRlseDone_33 <= 1'b0;
            end
            if(_zz_351[34]) begin
              rRlseDone_34 <= 1'b0;
            end
            if(_zz_351[35]) begin
              rRlseDone_35 <= 1'b0;
            end
            if(_zz_351[36]) begin
              rRlseDone_36 <= 1'b0;
            end
            if(_zz_351[37]) begin
              rRlseDone_37 <= 1'b0;
            end
            if(_zz_351[38]) begin
              rRlseDone_38 <= 1'b0;
            end
            if(_zz_351[39]) begin
              rRlseDone_39 <= 1'b0;
            end
            if(_zz_351[40]) begin
              rRlseDone_40 <= 1'b0;
            end
            if(_zz_351[41]) begin
              rRlseDone_41 <= 1'b0;
            end
            if(_zz_351[42]) begin
              rRlseDone_42 <= 1'b0;
            end
            if(_zz_351[43]) begin
              rRlseDone_43 <= 1'b0;
            end
            if(_zz_351[44]) begin
              rRlseDone_44 <= 1'b0;
            end
            if(_zz_351[45]) begin
              rRlseDone_45 <= 1'b0;
            end
            if(_zz_351[46]) begin
              rRlseDone_46 <= 1'b0;
            end
            if(_zz_351[47]) begin
              rRlseDone_47 <= 1'b0;
            end
            if(_zz_351[48]) begin
              rRlseDone_48 <= 1'b0;
            end
            if(_zz_351[49]) begin
              rRlseDone_49 <= 1'b0;
            end
            if(_zz_351[50]) begin
              rRlseDone_50 <= 1'b0;
            end
            if(_zz_351[51]) begin
              rRlseDone_51 <= 1'b0;
            end
            if(_zz_351[52]) begin
              rRlseDone_52 <= 1'b0;
            end
            if(_zz_351[53]) begin
              rRlseDone_53 <= 1'b0;
            end
            if(_zz_351[54]) begin
              rRlseDone_54 <= 1'b0;
            end
            if(_zz_351[55]) begin
              rRlseDone_55 <= 1'b0;
            end
            if(_zz_351[56]) begin
              rRlseDone_56 <= 1'b0;
            end
            if(_zz_351[57]) begin
              rRlseDone_57 <= 1'b0;
            end
            if(_zz_351[58]) begin
              rRlseDone_58 <= 1'b0;
            end
            if(_zz_351[59]) begin
              rRlseDone_59 <= 1'b0;
            end
            if(_zz_351[60]) begin
              rRlseDone_60 <= 1'b0;
            end
            if(_zz_351[61]) begin
              rRlseDone_61 <= 1'b0;
            end
            if(_zz_351[62]) begin
              rRlseDone_62 <= 1'b0;
            end
            if(_zz_351[63]) begin
              rRlseDone_63 <= 1'b0;
            end
            if(_zz_379[0]) begin
              rTimeOut_0 <= 1'b0;
            end
            if(_zz_379[1]) begin
              rTimeOut_1 <= 1'b0;
            end
            if(_zz_379[2]) begin
              rTimeOut_2 <= 1'b0;
            end
            if(_zz_379[3]) begin
              rTimeOut_3 <= 1'b0;
            end
            if(_zz_379[4]) begin
              rTimeOut_4 <= 1'b0;
            end
            if(_zz_379[5]) begin
              rTimeOut_5 <= 1'b0;
            end
            if(_zz_379[6]) begin
              rTimeOut_6 <= 1'b0;
            end
            if(_zz_379[7]) begin
              rTimeOut_7 <= 1'b0;
            end
            if(_zz_379[8]) begin
              rTimeOut_8 <= 1'b0;
            end
            if(_zz_379[9]) begin
              rTimeOut_9 <= 1'b0;
            end
            if(_zz_379[10]) begin
              rTimeOut_10 <= 1'b0;
            end
            if(_zz_379[11]) begin
              rTimeOut_11 <= 1'b0;
            end
            if(_zz_379[12]) begin
              rTimeOut_12 <= 1'b0;
            end
            if(_zz_379[13]) begin
              rTimeOut_13 <= 1'b0;
            end
            if(_zz_379[14]) begin
              rTimeOut_14 <= 1'b0;
            end
            if(_zz_379[15]) begin
              rTimeOut_15 <= 1'b0;
            end
            if(_zz_379[16]) begin
              rTimeOut_16 <= 1'b0;
            end
            if(_zz_379[17]) begin
              rTimeOut_17 <= 1'b0;
            end
            if(_zz_379[18]) begin
              rTimeOut_18 <= 1'b0;
            end
            if(_zz_379[19]) begin
              rTimeOut_19 <= 1'b0;
            end
            if(_zz_379[20]) begin
              rTimeOut_20 <= 1'b0;
            end
            if(_zz_379[21]) begin
              rTimeOut_21 <= 1'b0;
            end
            if(_zz_379[22]) begin
              rTimeOut_22 <= 1'b0;
            end
            if(_zz_379[23]) begin
              rTimeOut_23 <= 1'b0;
            end
            if(_zz_379[24]) begin
              rTimeOut_24 <= 1'b0;
            end
            if(_zz_379[25]) begin
              rTimeOut_25 <= 1'b0;
            end
            if(_zz_379[26]) begin
              rTimeOut_26 <= 1'b0;
            end
            if(_zz_379[27]) begin
              rTimeOut_27 <= 1'b0;
            end
            if(_zz_379[28]) begin
              rTimeOut_28 <= 1'b0;
            end
            if(_zz_379[29]) begin
              rTimeOut_29 <= 1'b0;
            end
            if(_zz_379[30]) begin
              rTimeOut_30 <= 1'b0;
            end
            if(_zz_379[31]) begin
              rTimeOut_31 <= 1'b0;
            end
            if(_zz_379[32]) begin
              rTimeOut_32 <= 1'b0;
            end
            if(_zz_379[33]) begin
              rTimeOut_33 <= 1'b0;
            end
            if(_zz_379[34]) begin
              rTimeOut_34 <= 1'b0;
            end
            if(_zz_379[35]) begin
              rTimeOut_35 <= 1'b0;
            end
            if(_zz_379[36]) begin
              rTimeOut_36 <= 1'b0;
            end
            if(_zz_379[37]) begin
              rTimeOut_37 <= 1'b0;
            end
            if(_zz_379[38]) begin
              rTimeOut_38 <= 1'b0;
            end
            if(_zz_379[39]) begin
              rTimeOut_39 <= 1'b0;
            end
            if(_zz_379[40]) begin
              rTimeOut_40 <= 1'b0;
            end
            if(_zz_379[41]) begin
              rTimeOut_41 <= 1'b0;
            end
            if(_zz_379[42]) begin
              rTimeOut_42 <= 1'b0;
            end
            if(_zz_379[43]) begin
              rTimeOut_43 <= 1'b0;
            end
            if(_zz_379[44]) begin
              rTimeOut_44 <= 1'b0;
            end
            if(_zz_379[45]) begin
              rTimeOut_45 <= 1'b0;
            end
            if(_zz_379[46]) begin
              rTimeOut_46 <= 1'b0;
            end
            if(_zz_379[47]) begin
              rTimeOut_47 <= 1'b0;
            end
            if(_zz_379[48]) begin
              rTimeOut_48 <= 1'b0;
            end
            if(_zz_379[49]) begin
              rTimeOut_49 <= 1'b0;
            end
            if(_zz_379[50]) begin
              rTimeOut_50 <= 1'b0;
            end
            if(_zz_379[51]) begin
              rTimeOut_51 <= 1'b0;
            end
            if(_zz_379[52]) begin
              rTimeOut_52 <= 1'b0;
            end
            if(_zz_379[53]) begin
              rTimeOut_53 <= 1'b0;
            end
            if(_zz_379[54]) begin
              rTimeOut_54 <= 1'b0;
            end
            if(_zz_379[55]) begin
              rTimeOut_55 <= 1'b0;
            end
            if(_zz_379[56]) begin
              rTimeOut_56 <= 1'b0;
            end
            if(_zz_379[57]) begin
              rTimeOut_57 <= 1'b0;
            end
            if(_zz_379[58]) begin
              rTimeOut_58 <= 1'b0;
            end
            if(_zz_379[59]) begin
              rTimeOut_59 <= 1'b0;
            end
            if(_zz_379[60]) begin
              rTimeOut_60 <= 1'b0;
            end
            if(_zz_379[61]) begin
              rTimeOut_61 <= 1'b0;
            end
            if(_zz_379[62]) begin
              rTimeOut_62 <= 1'b0;
            end
            if(_zz_379[63]) begin
              rTimeOut_63 <= 1'b0;
            end
            io_cntTxnLd <= (io_cntTxnLd + 32'h00000001);
            compLoadTxn_cntTxn <= (compLoadTxn_cntTxn + 32'h00000001);
          end
        end
        default : begin
        end
      endcase
      clkCnt_stateReg <= clkCnt_stateNext;
      case(clkCnt_stateReg)
        clkCnt_enumDef_IDLE : begin
          if(io_start) begin
            io_cntClk <= 32'h0;
            io_done <= 1'b0;
            io_cntTxnCmt <= 32'h0;
            io_cntTxnAbt <= 32'h0;
            io_cntTxnLd <= 32'h0;
            io_cntLockLoc <= 32'h0;
            io_cntLockRmt <= 32'h0;
            io_cntLockDenyLoc <= 32'h0;
            io_cntLockDenyRmt <= 32'h0;
          end
        end
        clkCnt_enumDef_CNT : begin
          io_cntClk <= (io_cntClk + 32'h00000001);
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(streamArbiter_8_io_output_ready) begin
      streamArbiter_8_io_output_rData_nId <= streamArbiter_8_io_output_payload_nId;
      streamArbiter_8_io_output_rData_tId <= streamArbiter_8_io_output_payload_tId;
      streamArbiter_8_io_output_rData_tabId <= streamArbiter_8_io_output_payload_tabId;
      streamArbiter_8_io_output_rData_snId <= streamArbiter_8_io_output_payload_snId;
      streamArbiter_8_io_output_rData_txnId <= streamArbiter_8_io_output_payload_txnId;
      streamArbiter_8_io_output_rData_lkType <= streamArbiter_8_io_output_payload_lkType;
      streamArbiter_8_io_output_rData_lkRelease <= streamArbiter_8_io_output_payload_lkRelease;
      streamArbiter_8_io_output_rData_txnTimeOut <= streamArbiter_8_io_output_payload_txnTimeOut;
      streamArbiter_8_io_output_rData_txnAbt <= streamArbiter_8_io_output_payload_txnAbt;
      streamArbiter_8_io_output_rData_lkIdx <= streamArbiter_8_io_output_payload_lkIdx;
      streamArbiter_8_io_output_rData_wLen <= streamArbiter_8_io_output_payload_wLen;
    end
    if(streamArbiter_8_io_output_s2mPipe_ready) begin
      streamArbiter_8_io_output_s2mPipe_rData_nId <= streamArbiter_8_io_output_s2mPipe_payload_nId;
      streamArbiter_8_io_output_s2mPipe_rData_tId <= streamArbiter_8_io_output_s2mPipe_payload_tId;
      streamArbiter_8_io_output_s2mPipe_rData_tabId <= streamArbiter_8_io_output_s2mPipe_payload_tabId;
      streamArbiter_8_io_output_s2mPipe_rData_snId <= streamArbiter_8_io_output_s2mPipe_payload_snId;
      streamArbiter_8_io_output_s2mPipe_rData_txnId <= streamArbiter_8_io_output_s2mPipe_payload_txnId;
      streamArbiter_8_io_output_s2mPipe_rData_lkType <= streamArbiter_8_io_output_s2mPipe_payload_lkType;
      streamArbiter_8_io_output_s2mPipe_rData_lkRelease <= streamArbiter_8_io_output_s2mPipe_payload_lkRelease;
      streamArbiter_8_io_output_s2mPipe_rData_txnTimeOut <= streamArbiter_8_io_output_s2mPipe_payload_txnTimeOut;
      streamArbiter_8_io_output_s2mPipe_rData_txnAbt <= streamArbiter_8_io_output_s2mPipe_payload_txnAbt;
      streamArbiter_8_io_output_s2mPipe_rData_lkIdx <= streamArbiter_8_io_output_s2mPipe_payload_lkIdx;
      streamArbiter_8_io_output_s2mPipe_rData_wLen <= streamArbiter_8_io_output_s2mPipe_payload_wLen;
    end
    if(streamArbiter_9_io_output_ready) begin
      streamArbiter_9_io_output_rData_nId <= streamArbiter_9_io_output_payload_nId;
      streamArbiter_9_io_output_rData_tId <= streamArbiter_9_io_output_payload_tId;
      streamArbiter_9_io_output_rData_tabId <= streamArbiter_9_io_output_payload_tabId;
      streamArbiter_9_io_output_rData_snId <= streamArbiter_9_io_output_payload_snId;
      streamArbiter_9_io_output_rData_txnId <= streamArbiter_9_io_output_payload_txnId;
      streamArbiter_9_io_output_rData_lkType <= streamArbiter_9_io_output_payload_lkType;
      streamArbiter_9_io_output_rData_lkRelease <= streamArbiter_9_io_output_payload_lkRelease;
      streamArbiter_9_io_output_rData_txnTimeOut <= streamArbiter_9_io_output_payload_txnTimeOut;
      streamArbiter_9_io_output_rData_txnAbt <= streamArbiter_9_io_output_payload_txnAbt;
      streamArbiter_9_io_output_rData_lkIdx <= streamArbiter_9_io_output_payload_lkIdx;
      streamArbiter_9_io_output_rData_wLen <= streamArbiter_9_io_output_payload_wLen;
    end
    if(streamArbiter_9_io_output_s2mPipe_ready) begin
      streamArbiter_9_io_output_s2mPipe_rData_nId <= streamArbiter_9_io_output_s2mPipe_payload_nId;
      streamArbiter_9_io_output_s2mPipe_rData_tId <= streamArbiter_9_io_output_s2mPipe_payload_tId;
      streamArbiter_9_io_output_s2mPipe_rData_tabId <= streamArbiter_9_io_output_s2mPipe_payload_tabId;
      streamArbiter_9_io_output_s2mPipe_rData_snId <= streamArbiter_9_io_output_s2mPipe_payload_snId;
      streamArbiter_9_io_output_s2mPipe_rData_txnId <= streamArbiter_9_io_output_s2mPipe_payload_txnId;
      streamArbiter_9_io_output_s2mPipe_rData_lkType <= streamArbiter_9_io_output_s2mPipe_payload_lkType;
      streamArbiter_9_io_output_s2mPipe_rData_lkRelease <= streamArbiter_9_io_output_s2mPipe_payload_lkRelease;
      streamArbiter_9_io_output_s2mPipe_rData_txnTimeOut <= streamArbiter_9_io_output_s2mPipe_payload_txnTimeOut;
      streamArbiter_9_io_output_s2mPipe_rData_txnAbt <= streamArbiter_9_io_output_s2mPipe_payload_txnAbt;
      streamArbiter_9_io_output_s2mPipe_rData_lkIdx <= streamArbiter_9_io_output_s2mPipe_payload_lkIdx;
      streamArbiter_9_io_output_s2mPipe_rData_wLen <= streamArbiter_9_io_output_s2mPipe_payload_wLen;
    end
    compLkReq_rIdxTxn2Start <= {_zz_compLkReq_rIdxTxn2Start_62,{_zz_compLkReq_rIdxTxn2Start_61,{_zz_compLkReq_rIdxTxn2Start_60,{_zz_compLkReq_rIdxTxn2Start_59,{_zz_compLkReq_rIdxTxn2Start_58,_zz_compLkReq_rIdxTxn2Start_57}}}}};
    if(io_lkRespLoc_fire) begin
      compLkRespLoc_rLkResp_valid <= io_lkRespLoc_valid;
      compLkRespLoc_rLkResp_ready <= io_lkRespLoc_ready;
      compLkRespLoc_rLkResp_payload_nId <= io_lkRespLoc_payload_nId;
      compLkRespLoc_rLkResp_payload_tId <= io_lkRespLoc_payload_tId;
      compLkRespLoc_rLkResp_payload_tabId <= io_lkRespLoc_payload_tabId;
      compLkRespLoc_rLkResp_payload_snId <= io_lkRespLoc_payload_snId;
      compLkRespLoc_rLkResp_payload_txnId <= io_lkRespLoc_payload_txnId;
      compLkRespLoc_rLkResp_payload_lkType <= io_lkRespLoc_payload_lkType;
      compLkRespLoc_rLkResp_payload_lkRelease <= io_lkRespLoc_payload_lkRelease;
      compLkRespLoc_rLkResp_payload_txnAbt <= io_lkRespLoc_payload_txnAbt;
      compLkRespLoc_rLkResp_payload_lkIdx <= io_lkRespLoc_payload_lkIdx;
      compLkRespLoc_rLkResp_payload_wLen <= io_lkRespLoc_payload_wLen;
      compLkRespLoc_rLkResp_payload_respType <= io_lkRespLoc_payload_respType;
      compLkRespLoc_rLkResp_payload_lkWaited <= io_lkRespLoc_payload_lkWaited;
    end
    if(io_lkRespLoc_fire_1) begin
      compLkRespLoc_rCurTxnId <= io_lkRespLoc_payload_txnId;
    end
    if(io_lkRespRmt_fire) begin
      compLkRespRmt_rLkResp_valid <= io_lkRespRmt_valid;
      compLkRespRmt_rLkResp_ready <= io_lkRespRmt_ready;
      compLkRespRmt_rLkResp_payload_nId <= io_lkRespRmt_payload_nId;
      compLkRespRmt_rLkResp_payload_tId <= io_lkRespRmt_payload_tId;
      compLkRespRmt_rLkResp_payload_tabId <= io_lkRespRmt_payload_tabId;
      compLkRespRmt_rLkResp_payload_snId <= io_lkRespRmt_payload_snId;
      compLkRespRmt_rLkResp_payload_txnId <= io_lkRespRmt_payload_txnId;
      compLkRespRmt_rLkResp_payload_lkType <= io_lkRespRmt_payload_lkType;
      compLkRespRmt_rLkResp_payload_lkRelease <= io_lkRespRmt_payload_lkRelease;
      compLkRespRmt_rLkResp_payload_txnAbt <= io_lkRespRmt_payload_txnAbt;
      compLkRespRmt_rLkResp_payload_lkIdx <= io_lkRespRmt_payload_lkIdx;
      compLkRespRmt_rLkResp_payload_wLen <= io_lkRespRmt_payload_wLen;
      compLkRespRmt_rLkResp_payload_respType <= io_lkRespRmt_payload_respType;
      compLkRespRmt_rLkResp_payload_lkWaited <= io_lkRespRmt_payload_lkWaited;
    end
    if(io_lkRespRmt_fire_1) begin
      compLkRespRmt_rCurTxnId <= io_lkRespRmt_payload_txnId;
    end
    compAxiResp_rAxiBFire <= io_axi_b_fire;
    compAxiResp_rAxiBId <= io_axi_b_payload_id;
    compTxnCmtLoc_rCmtTxn_nId <= compTxnCmtLoc_cmtTxn_nId;
    compTxnCmtLoc_rCmtTxn_tId <= compTxnCmtLoc_cmtTxn_tId;
    compTxnCmtLoc_rCmtTxn_tabId <= compTxnCmtLoc_cmtTxn_tabId;
    compTxnCmtLoc_rCmtTxn_lkType <= compTxnCmtLoc_cmtTxn_lkType;
    compTxnCmtLoc_rCmtTxn_wLen <= compTxnCmtLoc_cmtTxn_wLen;
    if(io_cmdAxi_r_fire) begin
      compLoadTxn_rCmdAxiData <= io_cmdAxi_r_payload_data;
    end
  end

  always @(posedge clk) begin
    _zz_81 <= (|compLkReq_mskTxn2Start);
  end


endmodule

module StreamFifo_2 (
  input               io_push_valid,
  output              io_push_ready,
  input      [511:0]  io_push_payload,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [511:0]  io_pop_payload,
  input               io_flush,
  output     [3:0]    io_occupancy,
  output     [3:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [511:0]  _zz_logic_ram_port0;
  wire       [2:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [2:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz_io_pop_payload;
  wire       [2:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [2:0]    logic_pushPtr_valueNext;
  reg        [2:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [2:0]    logic_popPtr_valueNext;
  reg        [2:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire                when_Stream_l1075;
  wire       [2:0]    logic_ptrDif;
  reg [511:0] logic_ram [0:7];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {2'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {2'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz_io_pop_payload = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_pop_payload) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= io_push_payload;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 3'b111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 3'b000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 3'b111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 3'b000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign io_pop_payload = _zz_logic_ram_port0;
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 3'b000;
      logic_popPtr_value <= 3'b000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1075) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamFifoLowLatency (
  input               io_push_valid,
  output              io_push_ready,
  input      [2:0]    io_push_payload,
  output reg          io_pop_valid,
  input               io_pop_ready,
  output reg [2:0]    io_pop_payload,
  input               io_flush,
  output     [3:0]    io_occupancy,
  input               clk,
  input               resetn
);

  wire       [2:0]    _zz_ram_port0;
  wire       [2:0]    _zz_pushPtr_valueNext;
  wire       [0:0]    _zz_pushPtr_valueNext_1;
  wire       [2:0]    _zz_popPtr_valueNext;
  wire       [0:0]    _zz_popPtr_valueNext_1;
  wire       [2:0]    _zz_ram_port;
  reg                 _zz_1;
  reg                 pushPtr_willIncrement;
  reg                 pushPtr_willClear;
  reg        [2:0]    pushPtr_valueNext;
  reg        [2:0]    pushPtr_value;
  wire                pushPtr_willOverflowIfInc;
  wire                pushPtr_willOverflow;
  reg                 popPtr_willIncrement;
  reg                 popPtr_willClear;
  reg        [2:0]    popPtr_valueNext;
  reg        [2:0]    popPtr_value;
  wire                popPtr_willOverflowIfInc;
  wire                popPtr_willOverflow;
  wire                ptrMatch;
  reg                 risingOccupancy;
  wire                empty;
  wire                full;
  wire                pushing;
  wire                popping;
  wire       [2:0]    readed;
  wire                when_Stream_l1175;
  wire                when_Stream_l1188;
  wire       [2:0]    ptrDif;
  (* ram_style = "distributed" *) reg [2:0] ram [0:7];

  assign _zz_pushPtr_valueNext_1 = pushPtr_willIncrement;
  assign _zz_pushPtr_valueNext = {2'd0, _zz_pushPtr_valueNext_1};
  assign _zz_popPtr_valueNext_1 = popPtr_willIncrement;
  assign _zz_popPtr_valueNext = {2'd0, _zz_popPtr_valueNext_1};
  assign _zz_ram_port = io_push_payload;
  assign _zz_ram_port0 = ram[popPtr_value];
  always @(posedge clk) begin
    if(_zz_1) begin
      ram[pushPtr_value] <= _zz_ram_port;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willIncrement = 1'b0;
    if(pushing) begin
      pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    pushPtr_willClear = 1'b0;
    if(io_flush) begin
      pushPtr_willClear = 1'b1;
    end
  end

  assign pushPtr_willOverflowIfInc = (pushPtr_value == 3'b111);
  assign pushPtr_willOverflow = (pushPtr_willOverflowIfInc && pushPtr_willIncrement);
  always @(*) begin
    pushPtr_valueNext = (pushPtr_value + _zz_pushPtr_valueNext);
    if(pushPtr_willClear) begin
      pushPtr_valueNext = 3'b000;
    end
  end

  always @(*) begin
    popPtr_willIncrement = 1'b0;
    if(popping) begin
      popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    popPtr_willClear = 1'b0;
    if(io_flush) begin
      popPtr_willClear = 1'b1;
    end
  end

  assign popPtr_willOverflowIfInc = (popPtr_value == 3'b111);
  assign popPtr_willOverflow = (popPtr_willOverflowIfInc && popPtr_willIncrement);
  always @(*) begin
    popPtr_valueNext = (popPtr_value + _zz_popPtr_valueNext);
    if(popPtr_willClear) begin
      popPtr_valueNext = 3'b000;
    end
  end

  assign ptrMatch = (pushPtr_value == popPtr_value);
  assign empty = (ptrMatch && (! risingOccupancy));
  assign full = (ptrMatch && risingOccupancy);
  assign pushing = (io_push_valid && io_push_ready);
  assign popping = (io_pop_valid && io_pop_ready);
  assign io_push_ready = (! full);
  assign readed = _zz_ram_port0;
  assign when_Stream_l1175 = (! empty);
  always @(*) begin
    if(when_Stream_l1175) begin
      io_pop_valid = 1'b1;
    end else begin
      io_pop_valid = io_push_valid;
    end
  end

  always @(*) begin
    if(when_Stream_l1175) begin
      io_pop_payload = readed;
    end else begin
      io_pop_payload = io_push_payload;
    end
  end

  assign when_Stream_l1188 = (pushing != popping);
  assign ptrDif = (pushPtr_value - popPtr_value);
  assign io_occupancy = {(risingOccupancy && ptrMatch),ptrDif};
  always @(posedge clk) begin
    if(!resetn) begin
      pushPtr_value <= 3'b000;
      popPtr_value <= 3'b000;
      risingOccupancy <= 1'b0;
    end else begin
      pushPtr_value <= pushPtr_valueNext;
      popPtr_value <= popPtr_valueNext;
      if(when_Stream_l1188) begin
        risingOccupancy <= pushing;
      end
      if(io_flush) begin
        risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

//StreamArbiter_2 replaced by StreamArbiter_2

//StreamDemux replaced by StreamDemux

//StreamFifo replaced by StreamFifo

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input      [0:0]    io_push_payload_nId,
  input      [21:0]   io_push_payload_tId,
  input      [2:0]    io_push_payload_tabId,
  input      [0:0]    io_push_payload_snId,
  input      [5:0]    io_push_payload_txnId,
  input      [1:0]    io_push_payload_lkType,
  input               io_push_payload_lkRelease,
  input               io_push_payload_txnTimeOut,
  input               io_push_payload_txnAbt,
  input      [5:0]    io_push_payload_lkIdx,
  input      [2:0]    io_push_payload_wLen,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [0:0]    io_pop_payload_nId,
  output     [21:0]   io_pop_payload_tId,
  output     [2:0]    io_pop_payload_tabId,
  output     [0:0]    io_pop_payload_snId,
  output     [5:0]    io_pop_payload_txnId,
  output     [1:0]    io_pop_payload_lkType,
  output              io_pop_payload_lkRelease,
  output              io_pop_payload_txnTimeOut,
  output              io_pop_payload_txnAbt,
  output     [5:0]    io_pop_payload_lkIdx,
  output     [2:0]    io_pop_payload_wLen,
  input               io_flush,
  output     [3:0]    io_occupancy,
  output     [3:0]    io_availability,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  reg        [46:0]   _zz_logic_ram_port0;
  wire       [2:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [2:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz__zz_io_pop_payload_nId;
  wire       [46:0]   _zz_logic_ram_port_1;
  wire       [2:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [2:0]    logic_pushPtr_valueNext;
  reg        [2:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [2:0]    logic_popPtr_valueNext;
  reg        [2:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire       [1:0]    _zz_io_pop_payload_lkType;
  wire       [46:0]   _zz_io_pop_payload_nId;
  wire       [1:0]    _zz_io_pop_payload_lkType_1;
  wire                when_Stream_l1075;
  wire       [2:0]    logic_ptrDif;
  `ifndef SYNTHESIS
  reg [47:0] io_push_payload_lkType_string;
  reg [47:0] io_pop_payload_lkType_string;
  reg [47:0] _zz_io_pop_payload_lkType_string;
  reg [47:0] _zz_io_pop_payload_lkType_1_string;
  `endif

  reg [46:0] logic_ram [0:7];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {2'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {2'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz__zz_io_pop_payload_nId = 1'b1;
  assign _zz_logic_ram_port_1 = {io_push_payload_wLen,{io_push_payload_lkIdx,{io_push_payload_txnAbt,{io_push_payload_txnTimeOut,{io_push_payload_lkRelease,{io_push_payload_lkType,{io_push_payload_txnId,{io_push_payload_snId,{io_push_payload_tabId,{io_push_payload_tId,io_push_payload_nId}}}}}}}}}};
  always @(posedge clk) begin
    if(_zz__zz_io_pop_payload_nId) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_push_payload_lkType)
      LkT_rd : io_push_payload_lkType_string = "rd    ";
      LkT_wr : io_push_payload_lkType_string = "wr    ";
      LkT_raw : io_push_payload_lkType_string = "raw   ";
      LkT_insTab : io_push_payload_lkType_string = "insTab";
      default : io_push_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_pop_payload_lkType)
      LkT_rd : io_pop_payload_lkType_string = "rd    ";
      LkT_wr : io_pop_payload_lkType_string = "wr    ";
      LkT_raw : io_pop_payload_lkType_string = "raw   ";
      LkT_insTab : io_pop_payload_lkType_string = "insTab";
      default : io_pop_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_pop_payload_lkType)
      LkT_rd : _zz_io_pop_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_pop_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_pop_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_pop_payload_lkType_string = "insTab";
      default : _zz_io_pop_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_pop_payload_lkType_1)
      LkT_rd : _zz_io_pop_payload_lkType_1_string = "rd    ";
      LkT_wr : _zz_io_pop_payload_lkType_1_string = "wr    ";
      LkT_raw : _zz_io_pop_payload_lkType_1_string = "raw   ";
      LkT_insTab : _zz_io_pop_payload_lkType_1_string = "insTab";
      default : _zz_io_pop_payload_lkType_1_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 3'b111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 3'b000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 3'b111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 3'b000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign _zz_io_pop_payload_nId = _zz_logic_ram_port0;
  assign _zz_io_pop_payload_lkType_1 = _zz_io_pop_payload_nId[34 : 33];
  assign _zz_io_pop_payload_lkType = _zz_io_pop_payload_lkType_1;
  assign io_pop_payload_nId = _zz_io_pop_payload_nId[0 : 0];
  assign io_pop_payload_tId = _zz_io_pop_payload_nId[22 : 1];
  assign io_pop_payload_tabId = _zz_io_pop_payload_nId[25 : 23];
  assign io_pop_payload_snId = _zz_io_pop_payload_nId[26 : 26];
  assign io_pop_payload_txnId = _zz_io_pop_payload_nId[32 : 27];
  assign io_pop_payload_lkType = _zz_io_pop_payload_lkType;
  assign io_pop_payload_lkRelease = _zz_io_pop_payload_nId[35];
  assign io_pop_payload_txnTimeOut = _zz_io_pop_payload_nId[36];
  assign io_pop_payload_txnAbt = _zz_io_pop_payload_nId[37];
  assign io_pop_payload_lkIdx = _zz_io_pop_payload_nId[43 : 38];
  assign io_pop_payload_wLen = _zz_io_pop_payload_nId[46 : 44];
  assign when_Stream_l1075 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 3'b000;
      logic_popPtr_value <= 3'b000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l1075) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamCrossbar_1 (
  input               io_inV_0_valid,
  output              io_inV_0_ready,
  input      [0:0]    io_inV_0_payload_nId,
  input      [21:0]   io_inV_0_payload_tId,
  input      [2:0]    io_inV_0_payload_tabId,
  input      [0:0]    io_inV_0_payload_snId,
  input      [5:0]    io_inV_0_payload_txnId,
  input      [1:0]    io_inV_0_payload_lkType,
  input               io_inV_0_payload_lkRelease,
  input               io_inV_0_payload_txnAbt,
  input      [5:0]    io_inV_0_payload_lkIdx,
  input      [2:0]    io_inV_0_payload_wLen,
  input      [1:0]    io_inV_0_payload_respType,
  input               io_inV_0_payload_lkWaited,
  output              io_outV_0_valid,
  input               io_outV_0_ready,
  output     [0:0]    io_outV_0_payload_nId,
  output     [21:0]   io_outV_0_payload_tId,
  output     [2:0]    io_outV_0_payload_tabId,
  output     [0:0]    io_outV_0_payload_snId,
  output     [5:0]    io_outV_0_payload_txnId,
  output     [1:0]    io_outV_0_payload_lkType,
  output              io_outV_0_payload_lkRelease,
  output              io_outV_0_payload_txnAbt,
  output     [5:0]    io_outV_0_payload_lkIdx,
  output     [2:0]    io_outV_0_payload_wLen,
  output     [1:0]    io_outV_0_payload_respType,
  output              io_outV_0_payload_lkWaited,
  output              io_outV_1_valid,
  input               io_outV_1_ready,
  output     [0:0]    io_outV_1_payload_nId,
  output     [21:0]   io_outV_1_payload_tId,
  output     [2:0]    io_outV_1_payload_tabId,
  output     [0:0]    io_outV_1_payload_snId,
  output     [5:0]    io_outV_1_payload_txnId,
  output     [1:0]    io_outV_1_payload_lkType,
  output              io_outV_1_payload_lkRelease,
  output              io_outV_1_payload_txnAbt,
  output     [5:0]    io_outV_1_payload_lkIdx,
  output     [2:0]    io_outV_1_payload_wLen,
  output     [1:0]    io_outV_1_payload_respType,
  output              io_outV_1_payload_lkWaited,
  input      [0:0]    io_inDemuxSel_0,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                inDemuxAry_0_io_outputs_0_ready;
  wire                inDemuxAry_0_io_outputs_1_ready;
  wire                inDemuxAry_0_io_input_ready;
  wire                inDemuxAry_0_io_outputs_0_valid;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_payload_respType;
  wire                inDemuxAry_0_io_outputs_0_payload_lkWaited;
  wire                inDemuxAry_0_io_outputs_1_valid;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_1_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_payload_lkType;
  wire                inDemuxAry_0_io_outputs_1_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_1_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_payload_respType;
  wire                inDemuxAry_0_io_outputs_1_payload_lkWaited;
  wire                outArbAry_0_io_inputs_0_ready;
  wire                outArbAry_0_io_output_valid;
  wire       [0:0]    outArbAry_0_io_output_payload_nId;
  wire       [21:0]   outArbAry_0_io_output_payload_tId;
  wire       [2:0]    outArbAry_0_io_output_payload_tabId;
  wire       [0:0]    outArbAry_0_io_output_payload_snId;
  wire       [5:0]    outArbAry_0_io_output_payload_txnId;
  wire       [1:0]    outArbAry_0_io_output_payload_lkType;
  wire                outArbAry_0_io_output_payload_lkRelease;
  wire                outArbAry_0_io_output_payload_txnAbt;
  wire       [5:0]    outArbAry_0_io_output_payload_lkIdx;
  wire       [2:0]    outArbAry_0_io_output_payload_wLen;
  wire       [1:0]    outArbAry_0_io_output_payload_respType;
  wire                outArbAry_0_io_output_payload_lkWaited;
  wire       [0:0]    outArbAry_0_io_chosenOH;
  wire                outArbAry_1_io_inputs_0_ready;
  wire                outArbAry_1_io_output_valid;
  wire       [0:0]    outArbAry_1_io_output_payload_nId;
  wire       [21:0]   outArbAry_1_io_output_payload_tId;
  wire       [2:0]    outArbAry_1_io_output_payload_tabId;
  wire       [0:0]    outArbAry_1_io_output_payload_snId;
  wire       [5:0]    outArbAry_1_io_output_payload_txnId;
  wire       [1:0]    outArbAry_1_io_output_payload_lkType;
  wire                outArbAry_1_io_output_payload_lkRelease;
  wire                outArbAry_1_io_output_payload_txnAbt;
  wire       [5:0]    outArbAry_1_io_output_payload_lkIdx;
  wire       [2:0]    outArbAry_1_io_output_payload_wLen;
  wire       [1:0]    outArbAry_1_io_output_payload_respType;
  wire                outArbAry_1_io_output_payload_lkWaited;
  wire       [0:0]    outArbAry_1_io_chosenOH;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_valid;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkWaited;
  reg                 inDemuxAry_0_io_outputs_0_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_0_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_0_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_0_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_rData_wLen;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_rData_respType;
  reg                 inDemuxAry_0_io_outputs_0_rData_lkWaited;
  wire       [1:0]    _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_valid;
  reg                 inDemuxAry_0_io_outputs_1_s2mPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_1_s2mPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkWaited;
  reg                 inDemuxAry_0_io_outputs_1_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_1_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_1_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_1_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_1_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_1_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_1_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_1_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_1_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_1_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_1_rData_wLen;
  reg        [1:0]    inDemuxAry_0_io_outputs_1_rData_respType;
  reg                 inDemuxAry_0_io_outputs_1_rData_lkWaited;
  wire       [1:0]    _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_valid;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType;
  wire                inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 inDemuxAry_0_io_outputs_1_s2mPipe_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_1_s2mPipe_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_wLen;
  reg        [1:0]    inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType;
  reg                 inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_1;
  `ifndef SYNTHESIS
  reg [47:0] io_inV_0_payload_lkType_string;
  reg [71:0] io_inV_0_payload_respType_string;
  reg [47:0] io_outV_0_payload_lkType_string;
  reg [71:0] io_outV_0_payload_respType_string;
  reg [47:0] io_outV_1_payload_lkType_string;
  reg [71:0] io_outV_1_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_rData_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_0_rData_respType_string;
  reg [47:0] _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_1_rData_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_1_rData_respType_string;
  reg [47:0] _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string;
  reg [71:0] inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string;
  `endif


  StreamDemux2_2 inDemuxAry_0 (
    .io_select                      (io_inDemuxSel_0                                ), //i
    .io_input_valid                 (io_inV_0_valid                                 ), //i
    .io_input_ready                 (inDemuxAry_0_io_input_ready                    ), //o
    .io_input_payload_nId           (io_inV_0_payload_nId                           ), //i
    .io_input_payload_tId           (io_inV_0_payload_tId[21:0]                     ), //i
    .io_input_payload_tabId         (io_inV_0_payload_tabId[2:0]                    ), //i
    .io_input_payload_snId          (io_inV_0_payload_snId                          ), //i
    .io_input_payload_txnId         (io_inV_0_payload_txnId[5:0]                    ), //i
    .io_input_payload_lkType        (io_inV_0_payload_lkType[1:0]                   ), //i
    .io_input_payload_lkRelease     (io_inV_0_payload_lkRelease                     ), //i
    .io_input_payload_txnAbt        (io_inV_0_payload_txnAbt                        ), //i
    .io_input_payload_lkIdx         (io_inV_0_payload_lkIdx[5:0]                    ), //i
    .io_input_payload_wLen          (io_inV_0_payload_wLen[2:0]                     ), //i
    .io_input_payload_respType      (io_inV_0_payload_respType[1:0]                 ), //i
    .io_input_payload_lkWaited      (io_inV_0_payload_lkWaited                      ), //i
    .io_outputs_0_valid             (inDemuxAry_0_io_outputs_0_valid                ), //o
    .io_outputs_0_ready             (inDemuxAry_0_io_outputs_0_ready                ), //i
    .io_outputs_0_payload_nId       (inDemuxAry_0_io_outputs_0_payload_nId          ), //o
    .io_outputs_0_payload_tId       (inDemuxAry_0_io_outputs_0_payload_tId[21:0]    ), //o
    .io_outputs_0_payload_tabId     (inDemuxAry_0_io_outputs_0_payload_tabId[2:0]   ), //o
    .io_outputs_0_payload_snId      (inDemuxAry_0_io_outputs_0_payload_snId         ), //o
    .io_outputs_0_payload_txnId     (inDemuxAry_0_io_outputs_0_payload_txnId[5:0]   ), //o
    .io_outputs_0_payload_lkType    (inDemuxAry_0_io_outputs_0_payload_lkType[1:0]  ), //o
    .io_outputs_0_payload_lkRelease (inDemuxAry_0_io_outputs_0_payload_lkRelease    ), //o
    .io_outputs_0_payload_txnAbt    (inDemuxAry_0_io_outputs_0_payload_txnAbt       ), //o
    .io_outputs_0_payload_lkIdx     (inDemuxAry_0_io_outputs_0_payload_lkIdx[5:0]   ), //o
    .io_outputs_0_payload_wLen      (inDemuxAry_0_io_outputs_0_payload_wLen[2:0]    ), //o
    .io_outputs_0_payload_respType  (inDemuxAry_0_io_outputs_0_payload_respType[1:0]), //o
    .io_outputs_0_payload_lkWaited  (inDemuxAry_0_io_outputs_0_payload_lkWaited     ), //o
    .io_outputs_1_valid             (inDemuxAry_0_io_outputs_1_valid                ), //o
    .io_outputs_1_ready             (inDemuxAry_0_io_outputs_1_ready                ), //i
    .io_outputs_1_payload_nId       (inDemuxAry_0_io_outputs_1_payload_nId          ), //o
    .io_outputs_1_payload_tId       (inDemuxAry_0_io_outputs_1_payload_tId[21:0]    ), //o
    .io_outputs_1_payload_tabId     (inDemuxAry_0_io_outputs_1_payload_tabId[2:0]   ), //o
    .io_outputs_1_payload_snId      (inDemuxAry_0_io_outputs_1_payload_snId         ), //o
    .io_outputs_1_payload_txnId     (inDemuxAry_0_io_outputs_1_payload_txnId[5:0]   ), //o
    .io_outputs_1_payload_lkType    (inDemuxAry_0_io_outputs_1_payload_lkType[1:0]  ), //o
    .io_outputs_1_payload_lkRelease (inDemuxAry_0_io_outputs_1_payload_lkRelease    ), //o
    .io_outputs_1_payload_txnAbt    (inDemuxAry_0_io_outputs_1_payload_txnAbt       ), //o
    .io_outputs_1_payload_lkIdx     (inDemuxAry_0_io_outputs_1_payload_lkIdx[5:0]   ), //o
    .io_outputs_1_payload_wLen      (inDemuxAry_0_io_outputs_1_payload_wLen[2:0]    ), //o
    .io_outputs_1_payload_respType  (inDemuxAry_0_io_outputs_1_payload_respType[1:0]), //o
    .io_outputs_1_payload_lkWaited  (inDemuxAry_0_io_outputs_1_payload_lkWaited     )  //o
  );
  StreamArbiter_3 outArbAry_0 (
    .io_inputs_0_valid             (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_0_ready             (outArbAry_0_io_inputs_0_ready                                  ), //o
    .io_inputs_0_payload_nId       (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_0_payload_tId       (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId[21:0]    ), //i
    .io_inputs_0_payload_tabId     (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_0_payload_snId      (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_0_payload_txnId     (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_0_payload_lkType    (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_0_payload_lkRelease (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_0_payload_txnAbt    (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_0_payload_lkIdx     (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_0_payload_wLen      (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_0_payload_respType  (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_0_payload_lkWaited  (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_output_valid               (outArbAry_0_io_output_valid                                    ), //o
    .io_output_ready               (io_outV_0_ready                                                ), //i
    .io_output_payload_nId         (outArbAry_0_io_output_payload_nId                              ), //o
    .io_output_payload_tId         (outArbAry_0_io_output_payload_tId[21:0]                        ), //o
    .io_output_payload_tabId       (outArbAry_0_io_output_payload_tabId[2:0]                       ), //o
    .io_output_payload_snId        (outArbAry_0_io_output_payload_snId                             ), //o
    .io_output_payload_txnId       (outArbAry_0_io_output_payload_txnId[5:0]                       ), //o
    .io_output_payload_lkType      (outArbAry_0_io_output_payload_lkType[1:0]                      ), //o
    .io_output_payload_lkRelease   (outArbAry_0_io_output_payload_lkRelease                        ), //o
    .io_output_payload_txnAbt      (outArbAry_0_io_output_payload_txnAbt                           ), //o
    .io_output_payload_lkIdx       (outArbAry_0_io_output_payload_lkIdx[5:0]                       ), //o
    .io_output_payload_wLen        (outArbAry_0_io_output_payload_wLen[2:0]                        ), //o
    .io_output_payload_respType    (outArbAry_0_io_output_payload_respType[1:0]                    ), //o
    .io_output_payload_lkWaited    (outArbAry_0_io_output_payload_lkWaited                         ), //o
    .io_chosenOH                   (outArbAry_0_io_chosenOH                                        ), //o
    .clk                           (clk                                                            ), //i
    .resetn                        (resetn                                                         )  //i
  );
  StreamArbiter_3 outArbAry_1 (
    .io_inputs_0_valid             (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_0_ready             (outArbAry_1_io_inputs_0_ready                                  ), //o
    .io_inputs_0_payload_nId       (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_0_payload_tId       (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tId[21:0]    ), //i
    .io_inputs_0_payload_tabId     (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_0_payload_snId      (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_0_payload_txnId     (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_0_payload_lkType    (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_0_payload_lkRelease (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_0_payload_txnAbt    (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_0_payload_lkIdx     (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_0_payload_wLen      (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_0_payload_respType  (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_0_payload_lkWaited  (inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_output_valid               (outArbAry_1_io_output_valid                                    ), //o
    .io_output_ready               (io_outV_1_ready                                                ), //i
    .io_output_payload_nId         (outArbAry_1_io_output_payload_nId                              ), //o
    .io_output_payload_tId         (outArbAry_1_io_output_payload_tId[21:0]                        ), //o
    .io_output_payload_tabId       (outArbAry_1_io_output_payload_tabId[2:0]                       ), //o
    .io_output_payload_snId        (outArbAry_1_io_output_payload_snId                             ), //o
    .io_output_payload_txnId       (outArbAry_1_io_output_payload_txnId[5:0]                       ), //o
    .io_output_payload_lkType      (outArbAry_1_io_output_payload_lkType[1:0]                      ), //o
    .io_output_payload_lkRelease   (outArbAry_1_io_output_payload_lkRelease                        ), //o
    .io_output_payload_txnAbt      (outArbAry_1_io_output_payload_txnAbt                           ), //o
    .io_output_payload_lkIdx       (outArbAry_1_io_output_payload_lkIdx[5:0]                       ), //o
    .io_output_payload_wLen        (outArbAry_1_io_output_payload_wLen[2:0]                        ), //o
    .io_output_payload_respType    (outArbAry_1_io_output_payload_respType[1:0]                    ), //o
    .io_output_payload_lkWaited    (outArbAry_1_io_output_payload_lkWaited                         ), //o
    .io_chosenOH                   (outArbAry_1_io_chosenOH                                        ), //o
    .clk                           (clk                                                            ), //i
    .resetn                        (resetn                                                         )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inV_0_payload_lkType)
      LkT_rd : io_inV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inV_0_payload_lkType_string = "insTab";
      default : io_inV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inV_0_payload_respType)
      LockRespType_grant : io_inV_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_inV_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inV_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inV_0_payload_respType_string = "release_1";
      default : io_inV_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_outV_0_payload_lkType)
      LkT_rd : io_outV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outV_0_payload_lkType_string = "insTab";
      default : io_outV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outV_0_payload_respType)
      LockRespType_grant : io_outV_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_outV_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_outV_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_outV_0_payload_respType_string = "release_1";
      default : io_outV_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_outV_1_payload_lkType)
      LkT_rd : io_outV_1_payload_lkType_string = "rd    ";
      LkT_wr : io_outV_1_payload_lkType_string = "wr    ";
      LkT_raw : io_outV_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_outV_1_payload_lkType_string = "insTab";
      default : io_outV_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outV_1_payload_respType)
      LockRespType_grant : io_outV_1_payload_respType_string = "grant    ";
      LockRespType_abort : io_outV_1_payload_respType_string = "abort    ";
      LockRespType_waiting : io_outV_1_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_outV_1_payload_respType_string = "release_1";
      default : io_outV_1_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_rData_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_0_rData_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_0_rData_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_0_rData_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_0_rData_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_0_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType)
      LockRespType_grant : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "release_1";
      default : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_1_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_1_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_1_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_1_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_1_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_rData_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_1_rData_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_1_rData_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_1_rData_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_1_rData_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_1_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType)
      LkT_rd : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType)
      LockRespType_grant : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "release_1";
      default : _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType)
      LockRespType_grant : inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string = "release_1";
      default : inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  `endif

  assign io_inV_0_ready = inDemuxAry_0_io_input_ready;
  assign inDemuxAry_0_io_outputs_0_ready = (! inDemuxAry_0_io_outputs_0_rValid);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_valid = (inDemuxAry_0_io_outputs_0_valid || inDemuxAry_0_io_outputs_0_rValid);
  assign _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkType : inDemuxAry_0_io_outputs_0_payload_lkType);
  assign _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_respType : inDemuxAry_0_io_outputs_0_payload_respType);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_nId : inDemuxAry_0_io_outputs_0_payload_nId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_tId : inDemuxAry_0_io_outputs_0_payload_tId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_tabId : inDemuxAry_0_io_outputs_0_payload_tabId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_snId : inDemuxAry_0_io_outputs_0_payload_snId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_txnId : inDemuxAry_0_io_outputs_0_payload_txnId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType = _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkRelease : inDemuxAry_0_io_outputs_0_payload_lkRelease);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_txnAbt : inDemuxAry_0_io_outputs_0_payload_txnAbt);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkIdx : inDemuxAry_0_io_outputs_0_payload_lkIdx);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_wLen : inDemuxAry_0_io_outputs_0_payload_wLen);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType = _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkWaited = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkWaited : inDemuxAry_0_io_outputs_0_payload_lkWaited);
  always @(*) begin
    inDemuxAry_0_io_outputs_0_s2mPipe_ready = inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      inDemuxAry_0_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid = inDemuxAry_0_io_outputs_0_s2mPipe_rValid;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt = inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen = inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_respType = inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkWaited = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkWaited;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready = outArbAry_0_io_inputs_0_ready;
  assign inDemuxAry_0_io_outputs_1_ready = (! inDemuxAry_0_io_outputs_1_rValid);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_valid = (inDemuxAry_0_io_outputs_1_valid || inDemuxAry_0_io_outputs_1_rValid);
  assign _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_lkType : inDemuxAry_0_io_outputs_1_payload_lkType);
  assign _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_respType : inDemuxAry_0_io_outputs_1_payload_respType);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_nId = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_nId : inDemuxAry_0_io_outputs_1_payload_nId);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_tId = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_tId : inDemuxAry_0_io_outputs_1_payload_tId);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_tabId = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_tabId : inDemuxAry_0_io_outputs_1_payload_tabId);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_snId = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_snId : inDemuxAry_0_io_outputs_1_payload_snId);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnId = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_txnId : inDemuxAry_0_io_outputs_1_payload_txnId);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType = _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkRelease = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_lkRelease : inDemuxAry_0_io_outputs_1_payload_lkRelease);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnAbt = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_txnAbt : inDemuxAry_0_io_outputs_1_payload_txnAbt);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkIdx = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_lkIdx : inDemuxAry_0_io_outputs_1_payload_lkIdx);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_wLen = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_wLen : inDemuxAry_0_io_outputs_1_payload_wLen);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType = _zz_inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkWaited = (inDemuxAry_0_io_outputs_1_rValid ? inDemuxAry_0_io_outputs_1_rData_lkWaited : inDemuxAry_0_io_outputs_1_payload_lkWaited);
  always @(*) begin
    inDemuxAry_0_io_outputs_1_s2mPipe_ready = inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      inDemuxAry_0_io_outputs_1_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_valid);
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_valid = inDemuxAry_0_io_outputs_1_s2mPipe_rValid;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_nId = inDemuxAry_0_io_outputs_1_s2mPipe_rData_nId;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tId = inDemuxAry_0_io_outputs_1_s2mPipe_rData_tId;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_tabId = inDemuxAry_0_io_outputs_1_s2mPipe_rData_tabId;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_snId = inDemuxAry_0_io_outputs_1_s2mPipe_rData_snId;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnId = inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnId;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkType = inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease = inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkRelease;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt = inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnAbt;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx = inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkIdx;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_wLen = inDemuxAry_0_io_outputs_1_s2mPipe_rData_wLen;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_respType = inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_payload_lkWaited = inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkWaited;
  assign inDemuxAry_0_io_outputs_1_s2mPipe_m2sPipe_ready = outArbAry_1_io_inputs_0_ready;
  assign io_outV_0_valid = outArbAry_0_io_output_valid;
  assign io_outV_0_payload_nId = outArbAry_0_io_output_payload_nId;
  assign io_outV_0_payload_tId = outArbAry_0_io_output_payload_tId;
  assign io_outV_0_payload_tabId = outArbAry_0_io_output_payload_tabId;
  assign io_outV_0_payload_snId = outArbAry_0_io_output_payload_snId;
  assign io_outV_0_payload_txnId = outArbAry_0_io_output_payload_txnId;
  assign io_outV_0_payload_lkType = outArbAry_0_io_output_payload_lkType;
  assign io_outV_0_payload_lkRelease = outArbAry_0_io_output_payload_lkRelease;
  assign io_outV_0_payload_txnAbt = outArbAry_0_io_output_payload_txnAbt;
  assign io_outV_0_payload_lkIdx = outArbAry_0_io_output_payload_lkIdx;
  assign io_outV_0_payload_wLen = outArbAry_0_io_output_payload_wLen;
  assign io_outV_0_payload_respType = outArbAry_0_io_output_payload_respType;
  assign io_outV_0_payload_lkWaited = outArbAry_0_io_output_payload_lkWaited;
  assign io_outV_1_valid = outArbAry_1_io_output_valid;
  assign io_outV_1_payload_nId = outArbAry_1_io_output_payload_nId;
  assign io_outV_1_payload_tId = outArbAry_1_io_output_payload_tId;
  assign io_outV_1_payload_tabId = outArbAry_1_io_output_payload_tabId;
  assign io_outV_1_payload_snId = outArbAry_1_io_output_payload_snId;
  assign io_outV_1_payload_txnId = outArbAry_1_io_output_payload_txnId;
  assign io_outV_1_payload_lkType = outArbAry_1_io_output_payload_lkType;
  assign io_outV_1_payload_lkRelease = outArbAry_1_io_output_payload_lkRelease;
  assign io_outV_1_payload_txnAbt = outArbAry_1_io_output_payload_txnAbt;
  assign io_outV_1_payload_lkIdx = outArbAry_1_io_output_payload_lkIdx;
  assign io_outV_1_payload_wLen = outArbAry_1_io_output_payload_wLen;
  assign io_outV_1_payload_respType = outArbAry_1_io_output_payload_respType;
  assign io_outV_1_payload_lkWaited = outArbAry_1_io_output_payload_lkWaited;
  always @(posedge clk) begin
    if(!resetn) begin
      inDemuxAry_0_io_outputs_0_rValid <= 1'b0;
      inDemuxAry_0_io_outputs_0_s2mPipe_rValid <= 1'b0;
      inDemuxAry_0_io_outputs_1_rValid <= 1'b0;
      inDemuxAry_0_io_outputs_1_s2mPipe_rValid <= 1'b0;
    end else begin
      if(inDemuxAry_0_io_outputs_0_valid) begin
        inDemuxAry_0_io_outputs_0_rValid <= 1'b1;
      end
      if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_0_rValid <= 1'b0;
      end
      if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_0_s2mPipe_rValid <= inDemuxAry_0_io_outputs_0_s2mPipe_valid;
      end
      if(inDemuxAry_0_io_outputs_1_valid) begin
        inDemuxAry_0_io_outputs_1_rValid <= 1'b1;
      end
      if(inDemuxAry_0_io_outputs_1_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_1_rValid <= 1'b0;
      end
      if(inDemuxAry_0_io_outputs_1_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_1_s2mPipe_rValid <= inDemuxAry_0_io_outputs_1_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(inDemuxAry_0_io_outputs_0_ready) begin
      inDemuxAry_0_io_outputs_0_rData_nId <= inDemuxAry_0_io_outputs_0_payload_nId;
      inDemuxAry_0_io_outputs_0_rData_tId <= inDemuxAry_0_io_outputs_0_payload_tId;
      inDemuxAry_0_io_outputs_0_rData_tabId <= inDemuxAry_0_io_outputs_0_payload_tabId;
      inDemuxAry_0_io_outputs_0_rData_snId <= inDemuxAry_0_io_outputs_0_payload_snId;
      inDemuxAry_0_io_outputs_0_rData_txnId <= inDemuxAry_0_io_outputs_0_payload_txnId;
      inDemuxAry_0_io_outputs_0_rData_lkType <= inDemuxAry_0_io_outputs_0_payload_lkType;
      inDemuxAry_0_io_outputs_0_rData_lkRelease <= inDemuxAry_0_io_outputs_0_payload_lkRelease;
      inDemuxAry_0_io_outputs_0_rData_txnAbt <= inDemuxAry_0_io_outputs_0_payload_txnAbt;
      inDemuxAry_0_io_outputs_0_rData_lkIdx <= inDemuxAry_0_io_outputs_0_payload_lkIdx;
      inDemuxAry_0_io_outputs_0_rData_wLen <= inDemuxAry_0_io_outputs_0_payload_wLen;
      inDemuxAry_0_io_outputs_0_rData_respType <= inDemuxAry_0_io_outputs_0_payload_respType;
      inDemuxAry_0_io_outputs_0_rData_lkWaited <= inDemuxAry_0_io_outputs_0_payload_lkWaited;
    end
    if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_respType <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_respType;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkWaited <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkWaited;
    end
    if(inDemuxAry_0_io_outputs_1_ready) begin
      inDemuxAry_0_io_outputs_1_rData_nId <= inDemuxAry_0_io_outputs_1_payload_nId;
      inDemuxAry_0_io_outputs_1_rData_tId <= inDemuxAry_0_io_outputs_1_payload_tId;
      inDemuxAry_0_io_outputs_1_rData_tabId <= inDemuxAry_0_io_outputs_1_payload_tabId;
      inDemuxAry_0_io_outputs_1_rData_snId <= inDemuxAry_0_io_outputs_1_payload_snId;
      inDemuxAry_0_io_outputs_1_rData_txnId <= inDemuxAry_0_io_outputs_1_payload_txnId;
      inDemuxAry_0_io_outputs_1_rData_lkType <= inDemuxAry_0_io_outputs_1_payload_lkType;
      inDemuxAry_0_io_outputs_1_rData_lkRelease <= inDemuxAry_0_io_outputs_1_payload_lkRelease;
      inDemuxAry_0_io_outputs_1_rData_txnAbt <= inDemuxAry_0_io_outputs_1_payload_txnAbt;
      inDemuxAry_0_io_outputs_1_rData_lkIdx <= inDemuxAry_0_io_outputs_1_payload_lkIdx;
      inDemuxAry_0_io_outputs_1_rData_wLen <= inDemuxAry_0_io_outputs_1_payload_wLen;
      inDemuxAry_0_io_outputs_1_rData_respType <= inDemuxAry_0_io_outputs_1_payload_respType;
      inDemuxAry_0_io_outputs_1_rData_lkWaited <= inDemuxAry_0_io_outputs_1_payload_lkWaited;
    end
    if(inDemuxAry_0_io_outputs_1_s2mPipe_ready) begin
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_nId <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_nId;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_tId <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_tId;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_tabId <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_tabId;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_snId <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_snId;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnId <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnId;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkType <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkType;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkRelease <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkRelease;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_txnAbt <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_txnAbt;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkIdx <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkIdx;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_wLen <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_wLen;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_respType <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_respType;
      inDemuxAry_0_io_outputs_1_s2mPipe_rData_lkWaited <= inDemuxAry_0_io_outputs_1_s2mPipe_payload_lkWaited;
    end
  end


endmodule

module StreamCrossbar (
  input               io_inV_0_valid,
  output              io_inV_0_ready,
  input      [0:0]    io_inV_0_payload_nId,
  input      [21:0]   io_inV_0_payload_tId,
  input      [2:0]    io_inV_0_payload_tabId,
  input      [0:0]    io_inV_0_payload_snId,
  input      [5:0]    io_inV_0_payload_txnId,
  input      [1:0]    io_inV_0_payload_lkType,
  input               io_inV_0_payload_lkRelease,
  input               io_inV_0_payload_txnTimeOut,
  input               io_inV_0_payload_txnAbt,
  input      [5:0]    io_inV_0_payload_lkIdx,
  input      [2:0]    io_inV_0_payload_wLen,
  input               io_inV_1_valid,
  output              io_inV_1_ready,
  input      [0:0]    io_inV_1_payload_nId,
  input      [21:0]   io_inV_1_payload_tId,
  input      [2:0]    io_inV_1_payload_tabId,
  input      [0:0]    io_inV_1_payload_snId,
  input      [5:0]    io_inV_1_payload_txnId,
  input      [1:0]    io_inV_1_payload_lkType,
  input               io_inV_1_payload_lkRelease,
  input               io_inV_1_payload_txnTimeOut,
  input               io_inV_1_payload_txnAbt,
  input      [5:0]    io_inV_1_payload_lkIdx,
  input      [2:0]    io_inV_1_payload_wLen,
  output              io_outV_0_valid,
  input               io_outV_0_ready,
  output     [0:0]    io_outV_0_payload_nId,
  output     [21:0]   io_outV_0_payload_tId,
  output     [2:0]    io_outV_0_payload_tabId,
  output     [0:0]    io_outV_0_payload_snId,
  output     [5:0]    io_outV_0_payload_txnId,
  output     [1:0]    io_outV_0_payload_lkType,
  output              io_outV_0_payload_lkRelease,
  output              io_outV_0_payload_txnTimeOut,
  output              io_outV_0_payload_txnAbt,
  output     [5:0]    io_outV_0_payload_lkIdx,
  output     [2:0]    io_outV_0_payload_wLen,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire                inDemuxAry_0_io_outputs_0_ready;
  wire                inDemuxAry_1_io_outputs_0_ready;
  wire                inDemuxAry_0_io_input_ready;
  wire                inDemuxAry_0_io_outputs_0_valid;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_payload_txnTimeOut;
  wire                inDemuxAry_0_io_outputs_0_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_payload_wLen;
  wire                inDemuxAry_1_io_input_ready;
  wire                inDemuxAry_1_io_outputs_0_valid;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_payload_nId;
  wire       [21:0]   inDemuxAry_1_io_outputs_0_payload_tId;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_payload_tabId;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_payload_snId;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_payload_txnId;
  wire       [1:0]    inDemuxAry_1_io_outputs_0_payload_lkType;
  wire                inDemuxAry_1_io_outputs_0_payload_lkRelease;
  wire                inDemuxAry_1_io_outputs_0_payload_txnTimeOut;
  wire                inDemuxAry_1_io_outputs_0_payload_txnAbt;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_payload_lkIdx;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_payload_wLen;
  wire                outArbAry_0_io_inputs_0_ready;
  wire                outArbAry_0_io_inputs_1_ready;
  wire                outArbAry_0_io_output_valid;
  wire       [0:0]    outArbAry_0_io_output_payload_nId;
  wire       [21:0]   outArbAry_0_io_output_payload_tId;
  wire       [2:0]    outArbAry_0_io_output_payload_tabId;
  wire       [0:0]    outArbAry_0_io_output_payload_snId;
  wire       [5:0]    outArbAry_0_io_output_payload_txnId;
  wire       [1:0]    outArbAry_0_io_output_payload_lkType;
  wire                outArbAry_0_io_output_payload_lkRelease;
  wire                outArbAry_0_io_output_payload_txnTimeOut;
  wire                outArbAry_0_io_output_payload_txnAbt;
  wire       [5:0]    outArbAry_0_io_output_payload_lkIdx;
  wire       [2:0]    outArbAry_0_io_output_payload_wLen;
  wire       [0:0]    outArbAry_0_io_chosen;
  wire       [1:0]    outArbAry_0_io_chosenOH;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_valid;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnTimeOut;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen;
  reg                 inDemuxAry_0_io_outputs_0_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_0_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_0_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_0_rData_txnTimeOut;
  reg                 inDemuxAry_0_io_outputs_0_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_rData_wLen;
  wire       [1:0]    _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rValid;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId;
  reg        [21:0]   inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId;
  reg        [0:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId;
  reg        [1:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnTimeOut;
  reg                 inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt;
  reg        [5:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx;
  reg        [2:0]    inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen;
  wire                when_Stream_l368;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_valid;
  reg                 inDemuxAry_1_io_outputs_0_s2mPipe_ready;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_nId;
  wire       [21:0]   inDemuxAry_1_io_outputs_0_s2mPipe_payload_tId;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_snId;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkRelease;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnTimeOut;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_payload_wLen;
  reg                 inDemuxAry_1_io_outputs_0_rValid;
  reg        [0:0]    inDemuxAry_1_io_outputs_0_rData_nId;
  reg        [21:0]   inDemuxAry_1_io_outputs_0_rData_tId;
  reg        [2:0]    inDemuxAry_1_io_outputs_0_rData_tabId;
  reg        [0:0]    inDemuxAry_1_io_outputs_0_rData_snId;
  reg        [5:0]    inDemuxAry_1_io_outputs_0_rData_txnId;
  reg        [1:0]    inDemuxAry_1_io_outputs_0_rData_lkType;
  reg                 inDemuxAry_1_io_outputs_0_rData_lkRelease;
  reg                 inDemuxAry_1_io_outputs_0_rData_txnTimeOut;
  reg                 inDemuxAry_1_io_outputs_0_rData_txnAbt;
  reg        [5:0]    inDemuxAry_1_io_outputs_0_rData_lkIdx;
  reg        [2:0]    inDemuxAry_1_io_outputs_0_rData_wLen;
  wire       [1:0]    _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_valid;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_ready;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_nId;
  wire       [21:0]   inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_wLen;
  reg                 inDemuxAry_1_io_outputs_0_s2mPipe_rValid;
  reg        [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_nId;
  reg        [21:0]   inDemuxAry_1_io_outputs_0_s2mPipe_rData_tId;
  reg        [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_tabId;
  reg        [0:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_snId;
  reg        [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnId;
  reg        [1:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType;
  reg                 inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkRelease;
  reg                 inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnTimeOut;
  reg                 inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnAbt;
  reg        [5:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkIdx;
  reg        [2:0]    inDemuxAry_1_io_outputs_0_s2mPipe_rData_wLen;
  wire                when_Stream_l368_1;
  `ifndef SYNTHESIS
  reg [47:0] io_inV_0_payload_lkType_string;
  reg [47:0] io_inV_1_payload_lkType_string;
  reg [47:0] io_outV_0_payload_lkType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_rData_lkType_string;
  reg [47:0] _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string;
  reg [47:0] inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_1_io_outputs_0_rData_lkType_string;
  reg [47:0] _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string;
  `endif


  StreamDemux2 inDemuxAry_0 (
    .io_input_valid                  (io_inV_0_valid                               ), //i
    .io_input_ready                  (inDemuxAry_0_io_input_ready                  ), //o
    .io_input_payload_nId            (io_inV_0_payload_nId                         ), //i
    .io_input_payload_tId            (io_inV_0_payload_tId[21:0]                   ), //i
    .io_input_payload_tabId          (io_inV_0_payload_tabId[2:0]                  ), //i
    .io_input_payload_snId           (io_inV_0_payload_snId                        ), //i
    .io_input_payload_txnId          (io_inV_0_payload_txnId[5:0]                  ), //i
    .io_input_payload_lkType         (io_inV_0_payload_lkType[1:0]                 ), //i
    .io_input_payload_lkRelease      (io_inV_0_payload_lkRelease                   ), //i
    .io_input_payload_txnTimeOut     (io_inV_0_payload_txnTimeOut                  ), //i
    .io_input_payload_txnAbt         (io_inV_0_payload_txnAbt                      ), //i
    .io_input_payload_lkIdx          (io_inV_0_payload_lkIdx[5:0]                  ), //i
    .io_input_payload_wLen           (io_inV_0_payload_wLen[2:0]                   ), //i
    .io_outputs_0_valid              (inDemuxAry_0_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (inDemuxAry_0_io_outputs_0_ready              ), //i
    .io_outputs_0_payload_nId        (inDemuxAry_0_io_outputs_0_payload_nId        ), //o
    .io_outputs_0_payload_tId        (inDemuxAry_0_io_outputs_0_payload_tId[21:0]  ), //o
    .io_outputs_0_payload_tabId      (inDemuxAry_0_io_outputs_0_payload_tabId[2:0] ), //o
    .io_outputs_0_payload_snId       (inDemuxAry_0_io_outputs_0_payload_snId       ), //o
    .io_outputs_0_payload_txnId      (inDemuxAry_0_io_outputs_0_payload_txnId[5:0] ), //o
    .io_outputs_0_payload_lkType     (inDemuxAry_0_io_outputs_0_payload_lkType[1:0]), //o
    .io_outputs_0_payload_lkRelease  (inDemuxAry_0_io_outputs_0_payload_lkRelease  ), //o
    .io_outputs_0_payload_txnTimeOut (inDemuxAry_0_io_outputs_0_payload_txnTimeOut ), //o
    .io_outputs_0_payload_txnAbt     (inDemuxAry_0_io_outputs_0_payload_txnAbt     ), //o
    .io_outputs_0_payload_lkIdx      (inDemuxAry_0_io_outputs_0_payload_lkIdx[5:0] ), //o
    .io_outputs_0_payload_wLen       (inDemuxAry_0_io_outputs_0_payload_wLen[2:0]  )  //o
  );
  StreamDemux2 inDemuxAry_1 (
    .io_input_valid                  (io_inV_1_valid                               ), //i
    .io_input_ready                  (inDemuxAry_1_io_input_ready                  ), //o
    .io_input_payload_nId            (io_inV_1_payload_nId                         ), //i
    .io_input_payload_tId            (io_inV_1_payload_tId[21:0]                   ), //i
    .io_input_payload_tabId          (io_inV_1_payload_tabId[2:0]                  ), //i
    .io_input_payload_snId           (io_inV_1_payload_snId                        ), //i
    .io_input_payload_txnId          (io_inV_1_payload_txnId[5:0]                  ), //i
    .io_input_payload_lkType         (io_inV_1_payload_lkType[1:0]                 ), //i
    .io_input_payload_lkRelease      (io_inV_1_payload_lkRelease                   ), //i
    .io_input_payload_txnTimeOut     (io_inV_1_payload_txnTimeOut                  ), //i
    .io_input_payload_txnAbt         (io_inV_1_payload_txnAbt                      ), //i
    .io_input_payload_lkIdx          (io_inV_1_payload_lkIdx[5:0]                  ), //i
    .io_input_payload_wLen           (io_inV_1_payload_wLen[2:0]                   ), //i
    .io_outputs_0_valid              (inDemuxAry_1_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (inDemuxAry_1_io_outputs_0_ready              ), //i
    .io_outputs_0_payload_nId        (inDemuxAry_1_io_outputs_0_payload_nId        ), //o
    .io_outputs_0_payload_tId        (inDemuxAry_1_io_outputs_0_payload_tId[21:0]  ), //o
    .io_outputs_0_payload_tabId      (inDemuxAry_1_io_outputs_0_payload_tabId[2:0] ), //o
    .io_outputs_0_payload_snId       (inDemuxAry_1_io_outputs_0_payload_snId       ), //o
    .io_outputs_0_payload_txnId      (inDemuxAry_1_io_outputs_0_payload_txnId[5:0] ), //o
    .io_outputs_0_payload_lkType     (inDemuxAry_1_io_outputs_0_payload_lkType[1:0]), //o
    .io_outputs_0_payload_lkRelease  (inDemuxAry_1_io_outputs_0_payload_lkRelease  ), //o
    .io_outputs_0_payload_txnTimeOut (inDemuxAry_1_io_outputs_0_payload_txnTimeOut ), //o
    .io_outputs_0_payload_txnAbt     (inDemuxAry_1_io_outputs_0_payload_txnAbt     ), //o
    .io_outputs_0_payload_lkIdx      (inDemuxAry_1_io_outputs_0_payload_lkIdx[5:0] ), //o
    .io_outputs_0_payload_wLen       (inDemuxAry_1_io_outputs_0_payload_wLen[2:0]  )  //o
  );
  StreamArbiter_2 outArbAry_0 (
    .io_inputs_0_valid              (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid              ), //i
    .io_inputs_0_ready              (outArbAry_0_io_inputs_0_ready                                ), //o
    .io_inputs_0_payload_nId        (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_inputs_0_payload_tId        (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId[21:0]  ), //i
    .io_inputs_0_payload_tabId      (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_inputs_0_payload_snId       (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_inputs_0_payload_txnId      (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_inputs_0_payload_lkType     (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_inputs_0_payload_lkRelease  (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_inputs_0_payload_txnTimeOut (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_inputs_0_payload_txnAbt     (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_inputs_0_payload_lkIdx      (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_inputs_0_payload_wLen       (inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_inputs_1_valid              (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_valid              ), //i
    .io_inputs_1_ready              (outArbAry_0_io_inputs_1_ready                                ), //o
    .io_inputs_1_payload_nId        (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_inputs_1_payload_tId        (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tId[21:0]  ), //i
    .io_inputs_1_payload_tabId      (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_inputs_1_payload_snId       (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_inputs_1_payload_txnId      (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_inputs_1_payload_lkType     (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_inputs_1_payload_lkRelease  (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_inputs_1_payload_txnTimeOut (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_inputs_1_payload_txnAbt     (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_inputs_1_payload_lkIdx      (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_inputs_1_payload_wLen       (inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_output_valid                (outArbAry_0_io_output_valid                                  ), //o
    .io_output_ready                (io_outV_0_ready                                              ), //i
    .io_output_payload_nId          (outArbAry_0_io_output_payload_nId                            ), //o
    .io_output_payload_tId          (outArbAry_0_io_output_payload_tId[21:0]                      ), //o
    .io_output_payload_tabId        (outArbAry_0_io_output_payload_tabId[2:0]                     ), //o
    .io_output_payload_snId         (outArbAry_0_io_output_payload_snId                           ), //o
    .io_output_payload_txnId        (outArbAry_0_io_output_payload_txnId[5:0]                     ), //o
    .io_output_payload_lkType       (outArbAry_0_io_output_payload_lkType[1:0]                    ), //o
    .io_output_payload_lkRelease    (outArbAry_0_io_output_payload_lkRelease                      ), //o
    .io_output_payload_txnTimeOut   (outArbAry_0_io_output_payload_txnTimeOut                     ), //o
    .io_output_payload_txnAbt       (outArbAry_0_io_output_payload_txnAbt                         ), //o
    .io_output_payload_lkIdx        (outArbAry_0_io_output_payload_lkIdx[5:0]                     ), //o
    .io_output_payload_wLen         (outArbAry_0_io_output_payload_wLen[2:0]                      ), //o
    .io_chosen                      (outArbAry_0_io_chosen                                        ), //o
    .io_chosenOH                    (outArbAry_0_io_chosenOH[1:0]                                 ), //o
    .clk                            (clk                                                          ), //i
    .resetn                         (resetn                                                       )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inV_0_payload_lkType)
      LkT_rd : io_inV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inV_0_payload_lkType_string = "insTab";
      default : io_inV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inV_1_payload_lkType)
      LkT_rd : io_inV_1_payload_lkType_string = "rd    ";
      LkT_wr : io_inV_1_payload_lkType_string = "wr    ";
      LkT_raw : io_inV_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_inV_1_payload_lkType_string = "insTab";
      default : io_inV_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outV_0_payload_lkType)
      LkT_rd : io_outV_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outV_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outV_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outV_0_payload_lkType_string = "insTab";
      default : io_outV_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType)
      LkT_rd : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "insTab";
      default : inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_1_io_outputs_0_rData_lkType)
      LkT_rd : inDemuxAry_1_io_outputs_0_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_1_io_outputs_0_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_1_io_outputs_0_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_1_io_outputs_0_rData_lkType_string = "insTab";
      default : inDemuxAry_1_io_outputs_0_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType)
      LkT_rd : inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string = "insTab";
      default : inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  `endif

  assign io_inV_0_ready = inDemuxAry_0_io_input_ready;
  assign io_inV_1_ready = inDemuxAry_1_io_input_ready;
  assign inDemuxAry_0_io_outputs_0_ready = (! inDemuxAry_0_io_outputs_0_rValid);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_valid = (inDemuxAry_0_io_outputs_0_valid || inDemuxAry_0_io_outputs_0_rValid);
  assign _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkType : inDemuxAry_0_io_outputs_0_payload_lkType);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_nId : inDemuxAry_0_io_outputs_0_payload_nId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_tId : inDemuxAry_0_io_outputs_0_payload_tId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_tabId : inDemuxAry_0_io_outputs_0_payload_tabId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_snId : inDemuxAry_0_io_outputs_0_payload_snId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_txnId : inDemuxAry_0_io_outputs_0_payload_txnId);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType = _zz_inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkRelease : inDemuxAry_0_io_outputs_0_payload_lkRelease);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnTimeOut = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_txnTimeOut : inDemuxAry_0_io_outputs_0_payload_txnTimeOut);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_txnAbt : inDemuxAry_0_io_outputs_0_payload_txnAbt);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_lkIdx : inDemuxAry_0_io_outputs_0_payload_lkIdx);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen = (inDemuxAry_0_io_outputs_0_rValid ? inDemuxAry_0_io_outputs_0_rData_wLen : inDemuxAry_0_io_outputs_0_payload_wLen);
  always @(*) begin
    inDemuxAry_0_io_outputs_0_s2mPipe_ready = inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      inDemuxAry_0_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid);
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_valid = inDemuxAry_0_io_outputs_0_s2mPipe_rValid;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_nId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_tabId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_snId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnId = inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkType = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut = inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnTimeOut;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt = inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx = inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_payload_wLen = inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen;
  assign inDemuxAry_0_io_outputs_0_s2mPipe_m2sPipe_ready = outArbAry_0_io_inputs_0_ready;
  assign inDemuxAry_1_io_outputs_0_ready = (! inDemuxAry_1_io_outputs_0_rValid);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_valid = (inDemuxAry_1_io_outputs_0_valid || inDemuxAry_1_io_outputs_0_rValid);
  assign _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_lkType : inDemuxAry_1_io_outputs_0_payload_lkType);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_nId = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_nId : inDemuxAry_1_io_outputs_0_payload_nId);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_tId = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_tId : inDemuxAry_1_io_outputs_0_payload_tId);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_tabId = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_tabId : inDemuxAry_1_io_outputs_0_payload_tabId);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_snId = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_snId : inDemuxAry_1_io_outputs_0_payload_snId);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnId = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_txnId : inDemuxAry_1_io_outputs_0_payload_txnId);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType = _zz_inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkRelease = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_lkRelease : inDemuxAry_1_io_outputs_0_payload_lkRelease);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnTimeOut = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_txnTimeOut : inDemuxAry_1_io_outputs_0_payload_txnTimeOut);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnAbt = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_txnAbt : inDemuxAry_1_io_outputs_0_payload_txnAbt);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkIdx = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_lkIdx : inDemuxAry_1_io_outputs_0_payload_lkIdx);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_payload_wLen = (inDemuxAry_1_io_outputs_0_rValid ? inDemuxAry_1_io_outputs_0_rData_wLen : inDemuxAry_1_io_outputs_0_payload_wLen);
  always @(*) begin
    inDemuxAry_1_io_outputs_0_s2mPipe_ready = inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      inDemuxAry_1_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_valid);
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_valid = inDemuxAry_1_io_outputs_0_s2mPipe_rValid;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_nId = inDemuxAry_1_io_outputs_0_s2mPipe_rData_nId;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tId = inDemuxAry_1_io_outputs_0_s2mPipe_rData_tId;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_tabId = inDemuxAry_1_io_outputs_0_s2mPipe_rData_tabId;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_snId = inDemuxAry_1_io_outputs_0_s2mPipe_rData_snId;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnId = inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnId;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkType = inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease = inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkRelease;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut = inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnTimeOut;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt = inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnAbt;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx = inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkIdx;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_payload_wLen = inDemuxAry_1_io_outputs_0_s2mPipe_rData_wLen;
  assign inDemuxAry_1_io_outputs_0_s2mPipe_m2sPipe_ready = outArbAry_0_io_inputs_1_ready;
  assign io_outV_0_valid = outArbAry_0_io_output_valid;
  assign io_outV_0_payload_nId = outArbAry_0_io_output_payload_nId;
  assign io_outV_0_payload_tId = outArbAry_0_io_output_payload_tId;
  assign io_outV_0_payload_tabId = outArbAry_0_io_output_payload_tabId;
  assign io_outV_0_payload_snId = outArbAry_0_io_output_payload_snId;
  assign io_outV_0_payload_txnId = outArbAry_0_io_output_payload_txnId;
  assign io_outV_0_payload_lkType = outArbAry_0_io_output_payload_lkType;
  assign io_outV_0_payload_lkRelease = outArbAry_0_io_output_payload_lkRelease;
  assign io_outV_0_payload_txnTimeOut = outArbAry_0_io_output_payload_txnTimeOut;
  assign io_outV_0_payload_txnAbt = outArbAry_0_io_output_payload_txnAbt;
  assign io_outV_0_payload_lkIdx = outArbAry_0_io_output_payload_lkIdx;
  assign io_outV_0_payload_wLen = outArbAry_0_io_output_payload_wLen;
  always @(posedge clk) begin
    if(!resetn) begin
      inDemuxAry_0_io_outputs_0_rValid <= 1'b0;
      inDemuxAry_0_io_outputs_0_s2mPipe_rValid <= 1'b0;
      inDemuxAry_1_io_outputs_0_rValid <= 1'b0;
      inDemuxAry_1_io_outputs_0_s2mPipe_rValid <= 1'b0;
    end else begin
      if(inDemuxAry_0_io_outputs_0_valid) begin
        inDemuxAry_0_io_outputs_0_rValid <= 1'b1;
      end
      if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_0_rValid <= 1'b0;
      end
      if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_0_io_outputs_0_s2mPipe_rValid <= inDemuxAry_0_io_outputs_0_s2mPipe_valid;
      end
      if(inDemuxAry_1_io_outputs_0_valid) begin
        inDemuxAry_1_io_outputs_0_rValid <= 1'b1;
      end
      if(inDemuxAry_1_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_1_io_outputs_0_rValid <= 1'b0;
      end
      if(inDemuxAry_1_io_outputs_0_s2mPipe_ready) begin
        inDemuxAry_1_io_outputs_0_s2mPipe_rValid <= inDemuxAry_1_io_outputs_0_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(inDemuxAry_0_io_outputs_0_ready) begin
      inDemuxAry_0_io_outputs_0_rData_nId <= inDemuxAry_0_io_outputs_0_payload_nId;
      inDemuxAry_0_io_outputs_0_rData_tId <= inDemuxAry_0_io_outputs_0_payload_tId;
      inDemuxAry_0_io_outputs_0_rData_tabId <= inDemuxAry_0_io_outputs_0_payload_tabId;
      inDemuxAry_0_io_outputs_0_rData_snId <= inDemuxAry_0_io_outputs_0_payload_snId;
      inDemuxAry_0_io_outputs_0_rData_txnId <= inDemuxAry_0_io_outputs_0_payload_txnId;
      inDemuxAry_0_io_outputs_0_rData_lkType <= inDemuxAry_0_io_outputs_0_payload_lkType;
      inDemuxAry_0_io_outputs_0_rData_lkRelease <= inDemuxAry_0_io_outputs_0_payload_lkRelease;
      inDemuxAry_0_io_outputs_0_rData_txnTimeOut <= inDemuxAry_0_io_outputs_0_payload_txnTimeOut;
      inDemuxAry_0_io_outputs_0_rData_txnAbt <= inDemuxAry_0_io_outputs_0_payload_txnAbt;
      inDemuxAry_0_io_outputs_0_rData_lkIdx <= inDemuxAry_0_io_outputs_0_payload_lkIdx;
      inDemuxAry_0_io_outputs_0_rData_wLen <= inDemuxAry_0_io_outputs_0_payload_wLen;
    end
    if(inDemuxAry_0_io_outputs_0_s2mPipe_ready) begin
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_nId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_nId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_tId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_tId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_tabId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_tabId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_snId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_snId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnId <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnId;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkType <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkType;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkRelease <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkRelease;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnTimeOut <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnTimeOut;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_txnAbt <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_txnAbt;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_lkIdx <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_lkIdx;
      inDemuxAry_0_io_outputs_0_s2mPipe_rData_wLen <= inDemuxAry_0_io_outputs_0_s2mPipe_payload_wLen;
    end
    if(inDemuxAry_1_io_outputs_0_ready) begin
      inDemuxAry_1_io_outputs_0_rData_nId <= inDemuxAry_1_io_outputs_0_payload_nId;
      inDemuxAry_1_io_outputs_0_rData_tId <= inDemuxAry_1_io_outputs_0_payload_tId;
      inDemuxAry_1_io_outputs_0_rData_tabId <= inDemuxAry_1_io_outputs_0_payload_tabId;
      inDemuxAry_1_io_outputs_0_rData_snId <= inDemuxAry_1_io_outputs_0_payload_snId;
      inDemuxAry_1_io_outputs_0_rData_txnId <= inDemuxAry_1_io_outputs_0_payload_txnId;
      inDemuxAry_1_io_outputs_0_rData_lkType <= inDemuxAry_1_io_outputs_0_payload_lkType;
      inDemuxAry_1_io_outputs_0_rData_lkRelease <= inDemuxAry_1_io_outputs_0_payload_lkRelease;
      inDemuxAry_1_io_outputs_0_rData_txnTimeOut <= inDemuxAry_1_io_outputs_0_payload_txnTimeOut;
      inDemuxAry_1_io_outputs_0_rData_txnAbt <= inDemuxAry_1_io_outputs_0_payload_txnAbt;
      inDemuxAry_1_io_outputs_0_rData_lkIdx <= inDemuxAry_1_io_outputs_0_payload_lkIdx;
      inDemuxAry_1_io_outputs_0_rData_wLen <= inDemuxAry_1_io_outputs_0_payload_wLen;
    end
    if(inDemuxAry_1_io_outputs_0_s2mPipe_ready) begin
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_nId <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_nId;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_tId <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_tId;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_tabId <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_tabId;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_snId <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_snId;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnId <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnId;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkType <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkType;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkRelease <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkRelease;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnTimeOut <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnTimeOut;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_txnAbt <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_txnAbt;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_lkIdx <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_lkIdx;
      inDemuxAry_1_io_outputs_0_s2mPipe_rData_wLen <= inDemuxAry_1_io_outputs_0_s2mPipe_payload_wLen;
    end
  end


endmodule

module LtCh (
  input               io_lkReq_valid,
  output              io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [21:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [21:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                ltAry_0_io_lkResp_ready;
  wire                ltAry_1_io_lkResp_ready;
  wire                ltAry_2_io_lkResp_ready;
  wire                ltAry_3_io_lkResp_ready;
  wire                ltAry_4_io_lkResp_ready;
  wire                ltAry_5_io_lkResp_ready;
  wire                ltAry_6_io_lkResp_ready;
  wire                ltAry_7_io_lkResp_ready;
  wire       [0:0]    streamDemux_7_io_select;
  wire       [2:0]    streamDemux_8_io_select;
  wire                streamDemux_8_io_outputs_0_ready;
  wire                streamDemux_8_io_outputs_1_ready;
  wire                streamDemux_8_io_outputs_2_ready;
  wire                streamDemux_8_io_outputs_3_ready;
  wire                streamDemux_8_io_outputs_4_ready;
  wire                streamDemux_8_io_outputs_5_ready;
  wire                streamDemux_8_io_outputs_6_ready;
  wire                streamDemux_8_io_outputs_7_ready;
  wire                ltAry_0_io_lkReq_ready;
  wire                ltAry_0_io_lkResp_valid;
  wire       [0:0]    ltAry_0_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_0_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_0_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_0_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_0_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_0_io_lkResp_payload_lkType;
  wire                ltAry_0_io_lkResp_payload_lkRelease;
  wire                ltAry_0_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_0_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_0_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_0_io_lkResp_payload_respType;
  wire                ltAry_0_io_lkResp_payload_lkWaited;
  wire                ltAry_1_io_lkReq_ready;
  wire                ltAry_1_io_lkResp_valid;
  wire       [0:0]    ltAry_1_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_1_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_1_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_1_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_1_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_1_io_lkResp_payload_lkType;
  wire                ltAry_1_io_lkResp_payload_lkRelease;
  wire                ltAry_1_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_1_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_1_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_1_io_lkResp_payload_respType;
  wire                ltAry_1_io_lkResp_payload_lkWaited;
  wire                ltAry_2_io_lkReq_ready;
  wire                ltAry_2_io_lkResp_valid;
  wire       [0:0]    ltAry_2_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_2_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_2_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_2_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_2_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_2_io_lkResp_payload_lkType;
  wire                ltAry_2_io_lkResp_payload_lkRelease;
  wire                ltAry_2_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_2_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_2_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_2_io_lkResp_payload_respType;
  wire                ltAry_2_io_lkResp_payload_lkWaited;
  wire                ltAry_3_io_lkReq_ready;
  wire                ltAry_3_io_lkResp_valid;
  wire       [0:0]    ltAry_3_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_3_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_3_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_3_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_3_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_3_io_lkResp_payload_lkType;
  wire                ltAry_3_io_lkResp_payload_lkRelease;
  wire                ltAry_3_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_3_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_3_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_3_io_lkResp_payload_respType;
  wire                ltAry_3_io_lkResp_payload_lkWaited;
  wire                ltAry_4_io_lkReq_ready;
  wire                ltAry_4_io_lkResp_valid;
  wire       [0:0]    ltAry_4_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_4_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_4_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_4_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_4_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_4_io_lkResp_payload_lkType;
  wire                ltAry_4_io_lkResp_payload_lkRelease;
  wire                ltAry_4_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_4_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_4_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_4_io_lkResp_payload_respType;
  wire                ltAry_4_io_lkResp_payload_lkWaited;
  wire                ltAry_5_io_lkReq_ready;
  wire                ltAry_5_io_lkResp_valid;
  wire       [0:0]    ltAry_5_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_5_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_5_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_5_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_5_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_5_io_lkResp_payload_lkType;
  wire                ltAry_5_io_lkResp_payload_lkRelease;
  wire                ltAry_5_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_5_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_5_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_5_io_lkResp_payload_respType;
  wire                ltAry_5_io_lkResp_payload_lkWaited;
  wire                ltAry_6_io_lkReq_ready;
  wire                ltAry_6_io_lkResp_valid;
  wire       [0:0]    ltAry_6_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_6_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_6_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_6_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_6_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_6_io_lkResp_payload_lkType;
  wire                ltAry_6_io_lkResp_payload_lkRelease;
  wire                ltAry_6_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_6_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_6_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_6_io_lkResp_payload_respType;
  wire                ltAry_6_io_lkResp_payload_lkWaited;
  wire                ltAry_7_io_lkReq_ready;
  wire                ltAry_7_io_lkResp_valid;
  wire       [0:0]    ltAry_7_io_lkResp_payload_nId;
  wire       [18:0]   ltAry_7_io_lkResp_payload_tId;
  wire       [2:0]    ltAry_7_io_lkResp_payload_tabId;
  wire       [0:0]    ltAry_7_io_lkResp_payload_snId;
  wire       [5:0]    ltAry_7_io_lkResp_payload_txnId;
  wire       [1:0]    ltAry_7_io_lkResp_payload_lkType;
  wire                ltAry_7_io_lkResp_payload_lkRelease;
  wire                ltAry_7_io_lkResp_payload_txnAbt;
  wire       [5:0]    ltAry_7_io_lkResp_payload_lkIdx;
  wire       [2:0]    ltAry_7_io_lkResp_payload_wLen;
  wire       [1:0]    ltAry_7_io_lkResp_payload_respType;
  wire                ltAry_7_io_lkResp_payload_lkWaited;
  wire                streamDemux_7_io_input_ready;
  wire                streamDemux_7_io_outputs_0_valid;
  wire       [0:0]    streamDemux_7_io_outputs_0_payload_nId;
  wire       [21:0]   streamDemux_7_io_outputs_0_payload_tId;
  wire       [2:0]    streamDemux_7_io_outputs_0_payload_tabId;
  wire       [0:0]    streamDemux_7_io_outputs_0_payload_snId;
  wire       [5:0]    streamDemux_7_io_outputs_0_payload_txnId;
  wire       [1:0]    streamDemux_7_io_outputs_0_payload_lkType;
  wire                streamDemux_7_io_outputs_0_payload_lkRelease;
  wire                streamDemux_7_io_outputs_0_payload_txnTimeOut;
  wire                streamDemux_7_io_outputs_0_payload_txnAbt;
  wire       [5:0]    streamDemux_7_io_outputs_0_payload_lkIdx;
  wire       [2:0]    streamDemux_7_io_outputs_0_payload_wLen;
  wire                streamDemux_7_io_outputs_1_valid;
  wire       [0:0]    streamDemux_7_io_outputs_1_payload_nId;
  wire       [21:0]   streamDemux_7_io_outputs_1_payload_tId;
  wire       [2:0]    streamDemux_7_io_outputs_1_payload_tabId;
  wire       [0:0]    streamDemux_7_io_outputs_1_payload_snId;
  wire       [5:0]    streamDemux_7_io_outputs_1_payload_txnId;
  wire       [1:0]    streamDemux_7_io_outputs_1_payload_lkType;
  wire                streamDemux_7_io_outputs_1_payload_lkRelease;
  wire                streamDemux_7_io_outputs_1_payload_txnTimeOut;
  wire                streamDemux_7_io_outputs_1_payload_txnAbt;
  wire       [5:0]    streamDemux_7_io_outputs_1_payload_lkIdx;
  wire       [2:0]    streamDemux_7_io_outputs_1_payload_wLen;
  wire                streamDemux_8_io_input_ready;
  wire                streamDemux_8_io_outputs_0_valid;
  wire       [0:0]    streamDemux_8_io_outputs_0_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_0_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_0_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_0_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_0_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_0_payload_lkType;
  wire                streamDemux_8_io_outputs_0_payload_lkRelease;
  wire                streamDemux_8_io_outputs_0_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_0_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_0_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_0_payload_wLen;
  wire                streamDemux_8_io_outputs_1_valid;
  wire       [0:0]    streamDemux_8_io_outputs_1_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_1_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_1_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_1_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_1_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_1_payload_lkType;
  wire                streamDemux_8_io_outputs_1_payload_lkRelease;
  wire                streamDemux_8_io_outputs_1_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_1_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_1_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_1_payload_wLen;
  wire                streamDemux_8_io_outputs_2_valid;
  wire       [0:0]    streamDemux_8_io_outputs_2_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_2_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_2_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_2_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_2_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_2_payload_lkType;
  wire                streamDemux_8_io_outputs_2_payload_lkRelease;
  wire                streamDemux_8_io_outputs_2_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_2_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_2_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_2_payload_wLen;
  wire                streamDemux_8_io_outputs_3_valid;
  wire       [0:0]    streamDemux_8_io_outputs_3_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_3_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_3_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_3_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_3_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_3_payload_lkType;
  wire                streamDemux_8_io_outputs_3_payload_lkRelease;
  wire                streamDemux_8_io_outputs_3_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_3_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_3_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_3_payload_wLen;
  wire                streamDemux_8_io_outputs_4_valid;
  wire       [0:0]    streamDemux_8_io_outputs_4_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_4_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_4_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_4_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_4_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_4_payload_lkType;
  wire                streamDemux_8_io_outputs_4_payload_lkRelease;
  wire                streamDemux_8_io_outputs_4_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_4_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_4_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_4_payload_wLen;
  wire                streamDemux_8_io_outputs_5_valid;
  wire       [0:0]    streamDemux_8_io_outputs_5_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_5_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_5_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_5_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_5_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_5_payload_lkType;
  wire                streamDemux_8_io_outputs_5_payload_lkRelease;
  wire                streamDemux_8_io_outputs_5_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_5_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_5_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_5_payload_wLen;
  wire                streamDemux_8_io_outputs_6_valid;
  wire       [0:0]    streamDemux_8_io_outputs_6_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_6_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_6_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_6_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_6_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_6_payload_lkType;
  wire                streamDemux_8_io_outputs_6_payload_lkRelease;
  wire                streamDemux_8_io_outputs_6_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_6_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_6_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_6_payload_wLen;
  wire                streamDemux_8_io_outputs_7_valid;
  wire       [0:0]    streamDemux_8_io_outputs_7_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_7_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_7_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_7_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_7_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_7_payload_lkType;
  wire                streamDemux_8_io_outputs_7_payload_lkRelease;
  wire                streamDemux_8_io_outputs_7_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_7_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_7_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_7_payload_wLen;
  wire                lkRespArb_io_inputs_0_ready;
  wire                lkRespArb_io_inputs_1_ready;
  wire                lkRespArb_io_inputs_2_ready;
  wire                lkRespArb_io_inputs_3_ready;
  wire                lkRespArb_io_inputs_4_ready;
  wire                lkRespArb_io_inputs_5_ready;
  wire                lkRespArb_io_inputs_6_ready;
  wire                lkRespArb_io_inputs_7_ready;
  wire                lkRespArb_io_output_valid;
  wire       [0:0]    lkRespArb_io_output_payload_nId;
  wire       [18:0]   lkRespArb_io_output_payload_tId;
  wire       [2:0]    lkRespArb_io_output_payload_tabId;
  wire       [0:0]    lkRespArb_io_output_payload_snId;
  wire       [5:0]    lkRespArb_io_output_payload_txnId;
  wire       [1:0]    lkRespArb_io_output_payload_lkType;
  wire                lkRespArb_io_output_payload_lkRelease;
  wire                lkRespArb_io_output_payload_txnAbt;
  wire       [5:0]    lkRespArb_io_output_payload_lkIdx;
  wire       [2:0]    lkRespArb_io_output_payload_wLen;
  wire       [1:0]    lkRespArb_io_output_payload_respType;
  wire                lkRespArb_io_output_payload_lkWaited;
  wire       [2:0]    lkRespArb_io_chosen;
  wire       [7:0]    lkRespArb_io_chosenOH;
  wire                streamArbiter_8_io_inputs_0_ready;
  wire                streamArbiter_8_io_inputs_1_ready;
  wire                streamArbiter_8_io_output_valid;
  wire       [0:0]    streamArbiter_8_io_output_payload_nId;
  wire       [21:0]   streamArbiter_8_io_output_payload_tId;
  wire       [2:0]    streamArbiter_8_io_output_payload_tabId;
  wire       [0:0]    streamArbiter_8_io_output_payload_snId;
  wire       [5:0]    streamArbiter_8_io_output_payload_txnId;
  wire       [1:0]    streamArbiter_8_io_output_payload_lkType;
  wire                streamArbiter_8_io_output_payload_lkRelease;
  wire                streamArbiter_8_io_output_payload_txnAbt;
  wire       [5:0]    streamArbiter_8_io_output_payload_lkIdx;
  wire       [2:0]    streamArbiter_8_io_output_payload_wLen;
  wire       [1:0]    streamArbiter_8_io_output_payload_respType;
  wire                streamArbiter_8_io_output_payload_lkWaited;
  wire       [0:0]    streamArbiter_8_io_chosen;
  wire       [1:0]    streamArbiter_8_io_chosenOH;
  reg        [21:0]   _zz_lkRespInsTab_payload_tId;
  reg        [21:0]   _zz__zz_tupPtr_0;
  wire       [15:0]   _zz_lkReq2Lt_payload_tId;
  reg        [21:0]   tupPtr_0;
  reg        [21:0]   tupPtr_1;
  reg        [21:0]   tupPtr_2;
  reg        [21:0]   tupPtr_3;
  reg        [21:0]   tupPtr_4;
  reg        [21:0]   tupPtr_5;
  reg        [21:0]   tupPtr_6;
  reg        [21:0]   tupPtr_7;
  wire                lkRespInsTab_valid;
  wire                lkRespInsTab_ready;
  wire       [0:0]    lkRespInsTab_payload_nId;
  reg        [21:0]   lkRespInsTab_payload_tId;
  wire       [2:0]    lkRespInsTab_payload_tabId;
  wire       [0:0]    lkRespInsTab_payload_snId;
  wire       [5:0]    lkRespInsTab_payload_txnId;
  wire       [1:0]    lkRespInsTab_payload_lkType;
  wire                lkRespInsTab_payload_lkRelease;
  wire                lkRespInsTab_payload_txnAbt;
  wire       [5:0]    lkRespInsTab_payload_lkIdx;
  wire       [2:0]    lkRespInsTab_payload_wLen;
  wire       [1:0]    lkRespInsTab_payload_respType;
  wire                lkRespInsTab_payload_lkWaited;
  wire                lkRespTup_valid;
  wire                lkRespTup_ready;
  wire       [0:0]    lkRespTup_payload_nId;
  wire       [21:0]   lkRespTup_payload_tId;
  wire       [2:0]    lkRespTup_payload_tabId;
  wire       [0:0]    lkRespTup_payload_snId;
  wire       [5:0]    lkRespTup_payload_txnId;
  wire       [1:0]    lkRespTup_payload_lkType;
  wire                lkRespTup_payload_lkRelease;
  wire                lkRespTup_payload_txnAbt;
  wire       [5:0]    lkRespTup_payload_lkIdx;
  wire       [2:0]    lkRespTup_payload_wLen;
  wire       [1:0]    lkRespTup_payload_respType;
  wire                lkRespTup_payload_lkWaited;
  wire                lkRespInsTab_fire;
  wire       [7:0]    _zz_1;
  wire       [21:0]   _zz_tupPtr_0;
  wire                lkReq2Lt_valid;
  wire                lkReq2Lt_ready;
  wire       [0:0]    lkReq2Lt_payload_nId;
  wire       [18:0]   lkReq2Lt_payload_tId;
  wire       [2:0]    lkReq2Lt_payload_tabId;
  wire       [0:0]    lkReq2Lt_payload_snId;
  wire       [5:0]    lkReq2Lt_payload_txnId;
  wire       [1:0]    lkReq2Lt_payload_lkType;
  wire                lkReq2Lt_payload_lkRelease;
  wire                lkReq2Lt_payload_txnTimeOut;
  wire                lkReq2Lt_payload_txnAbt;
  wire       [5:0]    lkReq2Lt_payload_lkIdx;
  wire       [2:0]    lkReq2Lt_payload_wLen;
  wire                streamDemux_8_io_outputs_0_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_0_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_0_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_0_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_0_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_0_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_0_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_0_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_0_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_0_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_0_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_0_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_0_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_0_rData_lkType;
  reg                 streamDemux_8_io_outputs_0_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_0_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_0_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_0_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_0_rData_wLen;
  wire       [1:0]    _zz_payload_lkType;
  wire                streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_0_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_0_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_0_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_0_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_0_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_0_s2mPipe_rData_wLen;
  wire                when_Stream_l368;
  wire                streamDemux_8_io_outputs_1_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_1_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_1_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_1_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_1_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_1_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_1_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_1_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_1_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_1_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_1_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_1_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_1_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_1_rData_lkType;
  reg                 streamDemux_8_io_outputs_1_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_1_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_1_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_1_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_1_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_1;
  wire                streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_1_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_1_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_1_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_1_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_1_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_1_s2mPipe_rData_wLen;
  wire                when_Stream_l368_1;
  wire                streamDemux_8_io_outputs_2_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_2_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_2_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_2_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_2_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_2_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_2_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_2_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_2_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_2_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_2_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_2_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_2_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_2_rData_lkType;
  reg                 streamDemux_8_io_outputs_2_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_2_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_2_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_2_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_2_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_2;
  wire                streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_2_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_2_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_2_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_2_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_2_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_2_s2mPipe_rData_wLen;
  wire                when_Stream_l368_2;
  wire                streamDemux_8_io_outputs_3_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_3_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_3_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_3_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_3_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_3_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_3_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_3_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_3_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_3_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_3_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_3_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_3_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_3_rData_lkType;
  reg                 streamDemux_8_io_outputs_3_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_3_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_3_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_3_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_3_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_3;
  wire                streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_3_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_3_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_3_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_3_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_3_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_3_s2mPipe_rData_wLen;
  wire                when_Stream_l368_3;
  wire                streamDemux_8_io_outputs_4_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_4_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_4_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_4_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_4_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_4_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_4_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_4_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_4_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_4_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_4_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_4_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_4_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_4_rData_lkType;
  reg                 streamDemux_8_io_outputs_4_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_4_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_4_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_4_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_4_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_4;
  wire                streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_4_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_4_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_4_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_4_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_4_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_4_s2mPipe_rData_wLen;
  wire                when_Stream_l368_4;
  wire                streamDemux_8_io_outputs_5_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_5_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_5_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_5_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_5_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_5_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_5_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_5_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_5_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_5_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_5_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_5_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_5_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_5_rData_lkType;
  reg                 streamDemux_8_io_outputs_5_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_5_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_5_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_5_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_5_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_5;
  wire                streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_5_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_5_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_5_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_5_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_5_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_5_s2mPipe_rData_wLen;
  wire                when_Stream_l368_5;
  wire                streamDemux_8_io_outputs_6_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_6_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_6_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_6_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_6_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_6_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_6_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_6_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_6_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_6_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_6_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_6_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_6_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_6_rData_lkType;
  reg                 streamDemux_8_io_outputs_6_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_6_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_6_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_6_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_6_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_6;
  wire                streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_6_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_6_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_6_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_6_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_6_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_6_s2mPipe_rData_wLen;
  wire                when_Stream_l368_6;
  wire                streamDemux_8_io_outputs_7_s2mPipe_valid;
  reg                 streamDemux_8_io_outputs_7_s2mPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_7_s2mPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_7_s2mPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_7_s2mPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_7_s2mPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_7_s2mPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_7_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_7_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_7_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_7_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_7_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_7_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_7_rData_lkType;
  reg                 streamDemux_8_io_outputs_7_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_7_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_7_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_7_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_7_rData_wLen;
  wire       [1:0]    _zz_payload_lkType_7;
  wire                streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_valid;
  wire                streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_ready;
  wire       [0:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType;
  wire                streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkRelease;
  wire                streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnTimeOut;
  wire                streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_wLen;
  reg                 streamDemux_8_io_outputs_7_s2mPipe_rValid;
  reg        [0:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_nId;
  reg        [18:0]   streamDemux_8_io_outputs_7_s2mPipe_rData_tId;
  reg        [2:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_tabId;
  reg        [0:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_snId;
  reg        [5:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_txnId;
  reg        [1:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_lkType;
  reg                 streamDemux_8_io_outputs_7_s2mPipe_rData_lkRelease;
  reg                 streamDemux_8_io_outputs_7_s2mPipe_rData_txnTimeOut;
  reg                 streamDemux_8_io_outputs_7_s2mPipe_rData_txnAbt;
  reg        [5:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_lkIdx;
  reg        [2:0]    streamDemux_8_io_outputs_7_s2mPipe_rData_wLen;
  wire                when_Stream_l368_7;
  wire                ltAry_0_io_lkResp_s2mPipe_valid;
  reg                 ltAry_0_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_0_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_0_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_0_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_0_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_0_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_0_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_0_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_0_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_0_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_0_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_0_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_0_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_0_io_lkResp_rValid;
  reg        [0:0]    ltAry_0_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_0_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_0_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_0_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_0_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_0_io_lkResp_rData_lkType;
  reg                 ltAry_0_io_lkResp_rData_lkRelease;
  reg                 ltAry_0_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_0_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_0_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_0_io_lkResp_rData_respType;
  reg                 ltAry_0_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_0_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_0_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_0_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_0_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_0_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_0_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_0_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_0_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_0_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_0_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_0_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_0_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_0_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_0_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_0_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_8;
  wire                ltAry_1_io_lkResp_s2mPipe_valid;
  reg                 ltAry_1_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_1_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_1_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_1_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_1_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_1_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_1_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_1_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_1_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_1_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_1_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_1_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_1_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_1_io_lkResp_rValid;
  reg        [0:0]    ltAry_1_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_1_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_1_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_1_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_1_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_1_io_lkResp_rData_lkType;
  reg                 ltAry_1_io_lkResp_rData_lkRelease;
  reg                 ltAry_1_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_1_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_1_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_1_io_lkResp_rData_respType;
  reg                 ltAry_1_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_1_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_1_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_1_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_1_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_1_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_1_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_1_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_1_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_1_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_1_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_1_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_1_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_1_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_1_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_1_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_9;
  wire                ltAry_2_io_lkResp_s2mPipe_valid;
  reg                 ltAry_2_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_2_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_2_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_2_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_2_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_2_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_2_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_2_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_2_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_2_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_2_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_2_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_2_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_2_io_lkResp_rValid;
  reg        [0:0]    ltAry_2_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_2_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_2_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_2_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_2_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_2_io_lkResp_rData_lkType;
  reg                 ltAry_2_io_lkResp_rData_lkRelease;
  reg                 ltAry_2_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_2_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_2_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_2_io_lkResp_rData_respType;
  reg                 ltAry_2_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_2_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_2_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_2_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_2_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_2_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_2_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_2_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_2_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_2_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_2_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_2_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_2_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_2_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_2_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_2_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_10;
  wire                ltAry_3_io_lkResp_s2mPipe_valid;
  reg                 ltAry_3_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_3_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_3_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_3_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_3_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_3_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_3_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_3_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_3_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_3_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_3_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_3_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_3_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_3_io_lkResp_rValid;
  reg        [0:0]    ltAry_3_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_3_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_3_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_3_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_3_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_3_io_lkResp_rData_lkType;
  reg                 ltAry_3_io_lkResp_rData_lkRelease;
  reg                 ltAry_3_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_3_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_3_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_3_io_lkResp_rData_respType;
  reg                 ltAry_3_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_3_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_3_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_3_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_3_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_3_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_3_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_3_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_3_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_3_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_3_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_3_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_3_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_3_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_3_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_3_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_11;
  wire                ltAry_4_io_lkResp_s2mPipe_valid;
  reg                 ltAry_4_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_4_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_4_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_4_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_4_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_4_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_4_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_4_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_4_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_4_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_4_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_4_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_4_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_4_io_lkResp_rValid;
  reg        [0:0]    ltAry_4_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_4_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_4_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_4_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_4_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_4_io_lkResp_rData_lkType;
  reg                 ltAry_4_io_lkResp_rData_lkRelease;
  reg                 ltAry_4_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_4_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_4_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_4_io_lkResp_rData_respType;
  reg                 ltAry_4_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_4_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_4_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_4_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_4_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_4_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_4_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_4_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_4_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_4_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_4_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_4_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_4_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_4_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_4_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_4_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_12;
  wire                ltAry_5_io_lkResp_s2mPipe_valid;
  reg                 ltAry_5_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_5_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_5_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_5_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_5_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_5_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_5_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_5_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_5_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_5_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_5_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_5_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_5_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_5_io_lkResp_rValid;
  reg        [0:0]    ltAry_5_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_5_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_5_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_5_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_5_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_5_io_lkResp_rData_lkType;
  reg                 ltAry_5_io_lkResp_rData_lkRelease;
  reg                 ltAry_5_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_5_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_5_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_5_io_lkResp_rData_respType;
  reg                 ltAry_5_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_5_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_5_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_5_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_5_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_5_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_5_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_5_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_5_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_5_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_5_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_5_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_5_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_5_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_5_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_5_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_13;
  wire                ltAry_6_io_lkResp_s2mPipe_valid;
  reg                 ltAry_6_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_6_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_6_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_6_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_6_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_6_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_6_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_6_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_6_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_6_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_6_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_6_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_6_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_6_io_lkResp_rValid;
  reg        [0:0]    ltAry_6_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_6_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_6_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_6_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_6_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_6_io_lkResp_rData_lkType;
  reg                 ltAry_6_io_lkResp_rData_lkRelease;
  reg                 ltAry_6_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_6_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_6_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_6_io_lkResp_rData_respType;
  reg                 ltAry_6_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_6_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_6_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_6_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_6_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_6_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_6_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_6_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_6_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_6_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_6_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_6_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_6_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_6_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_6_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_6_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_14;
  wire                ltAry_7_io_lkResp_s2mPipe_valid;
  reg                 ltAry_7_io_lkResp_s2mPipe_ready;
  wire       [0:0]    ltAry_7_io_lkResp_s2mPipe_payload_nId;
  wire       [18:0]   ltAry_7_io_lkResp_s2mPipe_payload_tId;
  wire       [2:0]    ltAry_7_io_lkResp_s2mPipe_payload_tabId;
  wire       [0:0]    ltAry_7_io_lkResp_s2mPipe_payload_snId;
  wire       [5:0]    ltAry_7_io_lkResp_s2mPipe_payload_txnId;
  wire       [1:0]    ltAry_7_io_lkResp_s2mPipe_payload_lkType;
  wire                ltAry_7_io_lkResp_s2mPipe_payload_lkRelease;
  wire                ltAry_7_io_lkResp_s2mPipe_payload_txnAbt;
  wire       [5:0]    ltAry_7_io_lkResp_s2mPipe_payload_lkIdx;
  wire       [2:0]    ltAry_7_io_lkResp_s2mPipe_payload_wLen;
  wire       [1:0]    ltAry_7_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_7_io_lkResp_s2mPipe_payload_lkWaited;
  reg                 ltAry_7_io_lkResp_rValid;
  reg        [0:0]    ltAry_7_io_lkResp_rData_nId;
  reg        [18:0]   ltAry_7_io_lkResp_rData_tId;
  reg        [2:0]    ltAry_7_io_lkResp_rData_tabId;
  reg        [0:0]    ltAry_7_io_lkResp_rData_snId;
  reg        [5:0]    ltAry_7_io_lkResp_rData_txnId;
  reg        [1:0]    ltAry_7_io_lkResp_rData_lkType;
  reg                 ltAry_7_io_lkResp_rData_lkRelease;
  reg                 ltAry_7_io_lkResp_rData_txnAbt;
  reg        [5:0]    ltAry_7_io_lkResp_rData_lkIdx;
  reg        [2:0]    ltAry_7_io_lkResp_rData_wLen;
  reg        [1:0]    ltAry_7_io_lkResp_rData_respType;
  reg                 ltAry_7_io_lkResp_rData_lkWaited;
  wire       [1:0]    _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType;
  wire       [1:0]    _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType;
  wire                ltAry_7_io_lkResp_s2mPipe_m2sPipe_valid;
  wire                ltAry_7_io_lkResp_s2mPipe_m2sPipe_ready;
  wire       [0:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_nId;
  wire       [18:0]   ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tId;
  wire       [2:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tabId;
  wire       [0:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_snId;
  wire       [5:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnId;
  wire       [1:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType;
  wire                ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease;
  wire                ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt;
  wire       [5:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx;
  wire       [2:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_wLen;
  wire       [1:0]    ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType;
  wire                ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited;
  reg                 ltAry_7_io_lkResp_s2mPipe_rValid;
  reg        [0:0]    ltAry_7_io_lkResp_s2mPipe_rData_nId;
  reg        [18:0]   ltAry_7_io_lkResp_s2mPipe_rData_tId;
  reg        [2:0]    ltAry_7_io_lkResp_s2mPipe_rData_tabId;
  reg        [0:0]    ltAry_7_io_lkResp_s2mPipe_rData_snId;
  reg        [5:0]    ltAry_7_io_lkResp_s2mPipe_rData_txnId;
  reg        [1:0]    ltAry_7_io_lkResp_s2mPipe_rData_lkType;
  reg                 ltAry_7_io_lkResp_s2mPipe_rData_lkRelease;
  reg                 ltAry_7_io_lkResp_s2mPipe_rData_txnAbt;
  reg        [5:0]    ltAry_7_io_lkResp_s2mPipe_rData_lkIdx;
  reg        [2:0]    ltAry_7_io_lkResp_s2mPipe_rData_wLen;
  reg        [1:0]    ltAry_7_io_lkResp_s2mPipe_rData_respType;
  reg                 ltAry_7_io_lkResp_s2mPipe_rData_lkWaited;
  wire                when_Stream_l368_15;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] lkRespInsTab_payload_lkType_string;
  reg [71:0] lkRespInsTab_payload_respType_string;
  reg [47:0] lkRespTup_payload_lkType_string;
  reg [71:0] lkRespTup_payload_respType_string;
  reg [47:0] lkReq2Lt_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_0_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_1_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_1_string;
  reg [47:0] streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_2_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_2_string;
  reg [47:0] streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_3_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_3_string;
  reg [47:0] streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_4_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_4_string;
  reg [47:0] streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_5_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_5_string;
  reg [47:0] streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_6_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_6_string;
  reg [47:0] streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_7_rData_lkType_string;
  reg [47:0] _zz_payload_lkType_7_string;
  reg [47:0] streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string;
  reg [47:0] streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string;
  reg [47:0] ltAry_0_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_0_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_0_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_0_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_0_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_0_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_1_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_1_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_1_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_1_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_1_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_1_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_2_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_2_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_2_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_2_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_2_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_2_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_3_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_3_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_3_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_3_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_3_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_3_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_4_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_4_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_4_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_4_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_4_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_4_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_5_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_5_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_5_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_5_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_5_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_5_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_6_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_6_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_6_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_6_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_6_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_6_io_lkResp_s2mPipe_rData_respType_string;
  reg [47:0] ltAry_7_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] ltAry_7_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_7_io_lkResp_rData_lkType_string;
  reg [71:0] ltAry_7_io_lkResp_rData_respType_string;
  reg [47:0] _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string;
  reg [71:0] _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string;
  reg [47:0] ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string;
  reg [71:0] ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string;
  reg [47:0] ltAry_7_io_lkResp_s2mPipe_rData_lkType_string;
  reg [71:0] ltAry_7_io_lkResp_s2mPipe_rData_respType_string;
  `endif


  assign _zz_lkReq2Lt_payload_tId = io_lkReq_payload_tId[18 : 3];
  LockTableBW ltAry_0 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_0_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_0_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_0_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_0_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_0_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_0_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_0_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_0_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_0_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_0_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_0_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_0_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_0_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_0_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_0_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_1 ltAry_1 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_1_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_1_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_1_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_1_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_1_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_1_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_1_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_1_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_1_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_1_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_1_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_1_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_1_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_1_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_1_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_2 ltAry_2 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_2_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_2_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_2_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_2_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_2_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_2_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_2_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_2_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_2_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_2_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_2_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_2_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_2_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_2_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_2_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_3 ltAry_3 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_3_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_3_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_3_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_3_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_3_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_3_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_3_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_3_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_3_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_3_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_3_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_3_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_3_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_3_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_3_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_4 ltAry_4 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_4_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_4_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_4_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_4_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_4_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_4_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_4_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_4_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_4_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_4_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_4_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_4_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_4_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_4_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_4_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_5 ltAry_5 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_5_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_5_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_5_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_5_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_5_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_5_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_5_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_5_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_5_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_5_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_5_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_5_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_5_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_5_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_5_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_6 ltAry_6 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_6_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_6_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_6_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_6_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_6_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_6_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_6_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_6_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_6_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_6_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_6_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_6_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_6_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_6_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_6_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  LockTableBW_7 ltAry_7 (
    .io_lkReq_valid              (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_valid              ), //i
    .io_lkReq_ready              (ltAry_7_io_lkReq_ready                                        ), //o
    .io_lkReq_payload_nId        (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_nId        ), //i
    .io_lkReq_payload_tId        (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tId[18:0]  ), //i
    .io_lkReq_payload_tabId      (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tabId[2:0] ), //i
    .io_lkReq_payload_snId       (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_snId       ), //i
    .io_lkReq_payload_txnId      (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnId[5:0] ), //i
    .io_lkReq_payload_lkType     (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType[1:0]), //i
    .io_lkReq_payload_lkRelease  (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkRelease  ), //i
    .io_lkReq_payload_txnTimeOut (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnTimeOut ), //i
    .io_lkReq_payload_txnAbt     (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnAbt     ), //i
    .io_lkReq_payload_lkIdx      (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkIdx[5:0] ), //i
    .io_lkReq_payload_wLen       (streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_wLen[2:0]  ), //i
    .io_lkResp_valid             (ltAry_7_io_lkResp_valid                                       ), //o
    .io_lkResp_ready             (ltAry_7_io_lkResp_ready                                       ), //i
    .io_lkResp_payload_nId       (ltAry_7_io_lkResp_payload_nId                                 ), //o
    .io_lkResp_payload_tId       (ltAry_7_io_lkResp_payload_tId[18:0]                           ), //o
    .io_lkResp_payload_tabId     (ltAry_7_io_lkResp_payload_tabId[2:0]                          ), //o
    .io_lkResp_payload_snId      (ltAry_7_io_lkResp_payload_snId                                ), //o
    .io_lkResp_payload_txnId     (ltAry_7_io_lkResp_payload_txnId[5:0]                          ), //o
    .io_lkResp_payload_lkType    (ltAry_7_io_lkResp_payload_lkType[1:0]                         ), //o
    .io_lkResp_payload_lkRelease (ltAry_7_io_lkResp_payload_lkRelease                           ), //o
    .io_lkResp_payload_txnAbt    (ltAry_7_io_lkResp_payload_txnAbt                              ), //o
    .io_lkResp_payload_lkIdx     (ltAry_7_io_lkResp_payload_lkIdx[5:0]                          ), //o
    .io_lkResp_payload_wLen      (ltAry_7_io_lkResp_payload_wLen[2:0]                           ), //o
    .io_lkResp_payload_respType  (ltAry_7_io_lkResp_payload_respType[1:0]                       ), //o
    .io_lkResp_payload_lkWaited  (ltAry_7_io_lkResp_payload_lkWaited                            ), //o
    .resetn                      (resetn                                                        ), //i
    .clk                         (clk                                                           )  //i
  );
  StreamDemux streamDemux_7 (
    .io_select                       (streamDemux_7_io_select                       ), //i
    .io_input_valid                  (io_lkReq_valid                                ), //i
    .io_input_ready                  (streamDemux_7_io_input_ready                  ), //o
    .io_input_payload_nId            (io_lkReq_payload_nId                          ), //i
    .io_input_payload_tId            (io_lkReq_payload_tId[21:0]                    ), //i
    .io_input_payload_tabId          (io_lkReq_payload_tabId[2:0]                   ), //i
    .io_input_payload_snId           (io_lkReq_payload_snId                         ), //i
    .io_input_payload_txnId          (io_lkReq_payload_txnId[5:0]                   ), //i
    .io_input_payload_lkType         (io_lkReq_payload_lkType[1:0]                  ), //i
    .io_input_payload_lkRelease      (io_lkReq_payload_lkRelease                    ), //i
    .io_input_payload_txnTimeOut     (io_lkReq_payload_txnTimeOut                   ), //i
    .io_input_payload_txnAbt         (io_lkReq_payload_txnAbt                       ), //i
    .io_input_payload_lkIdx          (io_lkReq_payload_lkIdx[5:0]                   ), //i
    .io_input_payload_wLen           (io_lkReq_payload_wLen[2:0]                    ), //i
    .io_outputs_0_valid              (streamDemux_7_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (lkReq2Lt_ready                                ), //i
    .io_outputs_0_payload_nId        (streamDemux_7_io_outputs_0_payload_nId        ), //o
    .io_outputs_0_payload_tId        (streamDemux_7_io_outputs_0_payload_tId[21:0]  ), //o
    .io_outputs_0_payload_tabId      (streamDemux_7_io_outputs_0_payload_tabId[2:0] ), //o
    .io_outputs_0_payload_snId       (streamDemux_7_io_outputs_0_payload_snId       ), //o
    .io_outputs_0_payload_txnId      (streamDemux_7_io_outputs_0_payload_txnId[5:0] ), //o
    .io_outputs_0_payload_lkType     (streamDemux_7_io_outputs_0_payload_lkType[1:0]), //o
    .io_outputs_0_payload_lkRelease  (streamDemux_7_io_outputs_0_payload_lkRelease  ), //o
    .io_outputs_0_payload_txnTimeOut (streamDemux_7_io_outputs_0_payload_txnTimeOut ), //o
    .io_outputs_0_payload_txnAbt     (streamDemux_7_io_outputs_0_payload_txnAbt     ), //o
    .io_outputs_0_payload_lkIdx      (streamDemux_7_io_outputs_0_payload_lkIdx[5:0] ), //o
    .io_outputs_0_payload_wLen       (streamDemux_7_io_outputs_0_payload_wLen[2:0]  ), //o
    .io_outputs_1_valid              (streamDemux_7_io_outputs_1_valid              ), //o
    .io_outputs_1_ready              (lkRespInsTab_ready                            ), //i
    .io_outputs_1_payload_nId        (streamDemux_7_io_outputs_1_payload_nId        ), //o
    .io_outputs_1_payload_tId        (streamDemux_7_io_outputs_1_payload_tId[21:0]  ), //o
    .io_outputs_1_payload_tabId      (streamDemux_7_io_outputs_1_payload_tabId[2:0] ), //o
    .io_outputs_1_payload_snId       (streamDemux_7_io_outputs_1_payload_snId       ), //o
    .io_outputs_1_payload_txnId      (streamDemux_7_io_outputs_1_payload_txnId[5:0] ), //o
    .io_outputs_1_payload_lkType     (streamDemux_7_io_outputs_1_payload_lkType[1:0]), //o
    .io_outputs_1_payload_lkRelease  (streamDemux_7_io_outputs_1_payload_lkRelease  ), //o
    .io_outputs_1_payload_txnTimeOut (streamDemux_7_io_outputs_1_payload_txnTimeOut ), //o
    .io_outputs_1_payload_txnAbt     (streamDemux_7_io_outputs_1_payload_txnAbt     ), //o
    .io_outputs_1_payload_lkIdx      (streamDemux_7_io_outputs_1_payload_lkIdx[5:0] ), //o
    .io_outputs_1_payload_wLen       (streamDemux_7_io_outputs_1_payload_wLen[2:0]  )  //o
  );
  StreamDemux_1 streamDemux_8 (
    .io_select                       (streamDemux_8_io_select[2:0]                  ), //i
    .io_input_valid                  (lkReq2Lt_valid                                ), //i
    .io_input_ready                  (streamDemux_8_io_input_ready                  ), //o
    .io_input_payload_nId            (lkReq2Lt_payload_nId                          ), //i
    .io_input_payload_tId            (lkReq2Lt_payload_tId[18:0]                    ), //i
    .io_input_payload_tabId          (lkReq2Lt_payload_tabId[2:0]                   ), //i
    .io_input_payload_snId           (lkReq2Lt_payload_snId                         ), //i
    .io_input_payload_txnId          (lkReq2Lt_payload_txnId[5:0]                   ), //i
    .io_input_payload_lkType         (lkReq2Lt_payload_lkType[1:0]                  ), //i
    .io_input_payload_lkRelease      (lkReq2Lt_payload_lkRelease                    ), //i
    .io_input_payload_txnTimeOut     (lkReq2Lt_payload_txnTimeOut                   ), //i
    .io_input_payload_txnAbt         (lkReq2Lt_payload_txnAbt                       ), //i
    .io_input_payload_lkIdx          (lkReq2Lt_payload_lkIdx[5:0]                   ), //i
    .io_input_payload_wLen           (lkReq2Lt_payload_wLen[2:0]                    ), //i
    .io_outputs_0_valid              (streamDemux_8_io_outputs_0_valid              ), //o
    .io_outputs_0_ready              (streamDemux_8_io_outputs_0_ready              ), //i
    .io_outputs_0_payload_nId        (streamDemux_8_io_outputs_0_payload_nId        ), //o
    .io_outputs_0_payload_tId        (streamDemux_8_io_outputs_0_payload_tId[18:0]  ), //o
    .io_outputs_0_payload_tabId      (streamDemux_8_io_outputs_0_payload_tabId[2:0] ), //o
    .io_outputs_0_payload_snId       (streamDemux_8_io_outputs_0_payload_snId       ), //o
    .io_outputs_0_payload_txnId      (streamDemux_8_io_outputs_0_payload_txnId[5:0] ), //o
    .io_outputs_0_payload_lkType     (streamDemux_8_io_outputs_0_payload_lkType[1:0]), //o
    .io_outputs_0_payload_lkRelease  (streamDemux_8_io_outputs_0_payload_lkRelease  ), //o
    .io_outputs_0_payload_txnTimeOut (streamDemux_8_io_outputs_0_payload_txnTimeOut ), //o
    .io_outputs_0_payload_txnAbt     (streamDemux_8_io_outputs_0_payload_txnAbt     ), //o
    .io_outputs_0_payload_lkIdx      (streamDemux_8_io_outputs_0_payload_lkIdx[5:0] ), //o
    .io_outputs_0_payload_wLen       (streamDemux_8_io_outputs_0_payload_wLen[2:0]  ), //o
    .io_outputs_1_valid              (streamDemux_8_io_outputs_1_valid              ), //o
    .io_outputs_1_ready              (streamDemux_8_io_outputs_1_ready              ), //i
    .io_outputs_1_payload_nId        (streamDemux_8_io_outputs_1_payload_nId        ), //o
    .io_outputs_1_payload_tId        (streamDemux_8_io_outputs_1_payload_tId[18:0]  ), //o
    .io_outputs_1_payload_tabId      (streamDemux_8_io_outputs_1_payload_tabId[2:0] ), //o
    .io_outputs_1_payload_snId       (streamDemux_8_io_outputs_1_payload_snId       ), //o
    .io_outputs_1_payload_txnId      (streamDemux_8_io_outputs_1_payload_txnId[5:0] ), //o
    .io_outputs_1_payload_lkType     (streamDemux_8_io_outputs_1_payload_lkType[1:0]), //o
    .io_outputs_1_payload_lkRelease  (streamDemux_8_io_outputs_1_payload_lkRelease  ), //o
    .io_outputs_1_payload_txnTimeOut (streamDemux_8_io_outputs_1_payload_txnTimeOut ), //o
    .io_outputs_1_payload_txnAbt     (streamDemux_8_io_outputs_1_payload_txnAbt     ), //o
    .io_outputs_1_payload_lkIdx      (streamDemux_8_io_outputs_1_payload_lkIdx[5:0] ), //o
    .io_outputs_1_payload_wLen       (streamDemux_8_io_outputs_1_payload_wLen[2:0]  ), //o
    .io_outputs_2_valid              (streamDemux_8_io_outputs_2_valid              ), //o
    .io_outputs_2_ready              (streamDemux_8_io_outputs_2_ready              ), //i
    .io_outputs_2_payload_nId        (streamDemux_8_io_outputs_2_payload_nId        ), //o
    .io_outputs_2_payload_tId        (streamDemux_8_io_outputs_2_payload_tId[18:0]  ), //o
    .io_outputs_2_payload_tabId      (streamDemux_8_io_outputs_2_payload_tabId[2:0] ), //o
    .io_outputs_2_payload_snId       (streamDemux_8_io_outputs_2_payload_snId       ), //o
    .io_outputs_2_payload_txnId      (streamDemux_8_io_outputs_2_payload_txnId[5:0] ), //o
    .io_outputs_2_payload_lkType     (streamDemux_8_io_outputs_2_payload_lkType[1:0]), //o
    .io_outputs_2_payload_lkRelease  (streamDemux_8_io_outputs_2_payload_lkRelease  ), //o
    .io_outputs_2_payload_txnTimeOut (streamDemux_8_io_outputs_2_payload_txnTimeOut ), //o
    .io_outputs_2_payload_txnAbt     (streamDemux_8_io_outputs_2_payload_txnAbt     ), //o
    .io_outputs_2_payload_lkIdx      (streamDemux_8_io_outputs_2_payload_lkIdx[5:0] ), //o
    .io_outputs_2_payload_wLen       (streamDemux_8_io_outputs_2_payload_wLen[2:0]  ), //o
    .io_outputs_3_valid              (streamDemux_8_io_outputs_3_valid              ), //o
    .io_outputs_3_ready              (streamDemux_8_io_outputs_3_ready              ), //i
    .io_outputs_3_payload_nId        (streamDemux_8_io_outputs_3_payload_nId        ), //o
    .io_outputs_3_payload_tId        (streamDemux_8_io_outputs_3_payload_tId[18:0]  ), //o
    .io_outputs_3_payload_tabId      (streamDemux_8_io_outputs_3_payload_tabId[2:0] ), //o
    .io_outputs_3_payload_snId       (streamDemux_8_io_outputs_3_payload_snId       ), //o
    .io_outputs_3_payload_txnId      (streamDemux_8_io_outputs_3_payload_txnId[5:0] ), //o
    .io_outputs_3_payload_lkType     (streamDemux_8_io_outputs_3_payload_lkType[1:0]), //o
    .io_outputs_3_payload_lkRelease  (streamDemux_8_io_outputs_3_payload_lkRelease  ), //o
    .io_outputs_3_payload_txnTimeOut (streamDemux_8_io_outputs_3_payload_txnTimeOut ), //o
    .io_outputs_3_payload_txnAbt     (streamDemux_8_io_outputs_3_payload_txnAbt     ), //o
    .io_outputs_3_payload_lkIdx      (streamDemux_8_io_outputs_3_payload_lkIdx[5:0] ), //o
    .io_outputs_3_payload_wLen       (streamDemux_8_io_outputs_3_payload_wLen[2:0]  ), //o
    .io_outputs_4_valid              (streamDemux_8_io_outputs_4_valid              ), //o
    .io_outputs_4_ready              (streamDemux_8_io_outputs_4_ready              ), //i
    .io_outputs_4_payload_nId        (streamDemux_8_io_outputs_4_payload_nId        ), //o
    .io_outputs_4_payload_tId        (streamDemux_8_io_outputs_4_payload_tId[18:0]  ), //o
    .io_outputs_4_payload_tabId      (streamDemux_8_io_outputs_4_payload_tabId[2:0] ), //o
    .io_outputs_4_payload_snId       (streamDemux_8_io_outputs_4_payload_snId       ), //o
    .io_outputs_4_payload_txnId      (streamDemux_8_io_outputs_4_payload_txnId[5:0] ), //o
    .io_outputs_4_payload_lkType     (streamDemux_8_io_outputs_4_payload_lkType[1:0]), //o
    .io_outputs_4_payload_lkRelease  (streamDemux_8_io_outputs_4_payload_lkRelease  ), //o
    .io_outputs_4_payload_txnTimeOut (streamDemux_8_io_outputs_4_payload_txnTimeOut ), //o
    .io_outputs_4_payload_txnAbt     (streamDemux_8_io_outputs_4_payload_txnAbt     ), //o
    .io_outputs_4_payload_lkIdx      (streamDemux_8_io_outputs_4_payload_lkIdx[5:0] ), //o
    .io_outputs_4_payload_wLen       (streamDemux_8_io_outputs_4_payload_wLen[2:0]  ), //o
    .io_outputs_5_valid              (streamDemux_8_io_outputs_5_valid              ), //o
    .io_outputs_5_ready              (streamDemux_8_io_outputs_5_ready              ), //i
    .io_outputs_5_payload_nId        (streamDemux_8_io_outputs_5_payload_nId        ), //o
    .io_outputs_5_payload_tId        (streamDemux_8_io_outputs_5_payload_tId[18:0]  ), //o
    .io_outputs_5_payload_tabId      (streamDemux_8_io_outputs_5_payload_tabId[2:0] ), //o
    .io_outputs_5_payload_snId       (streamDemux_8_io_outputs_5_payload_snId       ), //o
    .io_outputs_5_payload_txnId      (streamDemux_8_io_outputs_5_payload_txnId[5:0] ), //o
    .io_outputs_5_payload_lkType     (streamDemux_8_io_outputs_5_payload_lkType[1:0]), //o
    .io_outputs_5_payload_lkRelease  (streamDemux_8_io_outputs_5_payload_lkRelease  ), //o
    .io_outputs_5_payload_txnTimeOut (streamDemux_8_io_outputs_5_payload_txnTimeOut ), //o
    .io_outputs_5_payload_txnAbt     (streamDemux_8_io_outputs_5_payload_txnAbt     ), //o
    .io_outputs_5_payload_lkIdx      (streamDemux_8_io_outputs_5_payload_lkIdx[5:0] ), //o
    .io_outputs_5_payload_wLen       (streamDemux_8_io_outputs_5_payload_wLen[2:0]  ), //o
    .io_outputs_6_valid              (streamDemux_8_io_outputs_6_valid              ), //o
    .io_outputs_6_ready              (streamDemux_8_io_outputs_6_ready              ), //i
    .io_outputs_6_payload_nId        (streamDemux_8_io_outputs_6_payload_nId        ), //o
    .io_outputs_6_payload_tId        (streamDemux_8_io_outputs_6_payload_tId[18:0]  ), //o
    .io_outputs_6_payload_tabId      (streamDemux_8_io_outputs_6_payload_tabId[2:0] ), //o
    .io_outputs_6_payload_snId       (streamDemux_8_io_outputs_6_payload_snId       ), //o
    .io_outputs_6_payload_txnId      (streamDemux_8_io_outputs_6_payload_txnId[5:0] ), //o
    .io_outputs_6_payload_lkType     (streamDemux_8_io_outputs_6_payload_lkType[1:0]), //o
    .io_outputs_6_payload_lkRelease  (streamDemux_8_io_outputs_6_payload_lkRelease  ), //o
    .io_outputs_6_payload_txnTimeOut (streamDemux_8_io_outputs_6_payload_txnTimeOut ), //o
    .io_outputs_6_payload_txnAbt     (streamDemux_8_io_outputs_6_payload_txnAbt     ), //o
    .io_outputs_6_payload_lkIdx      (streamDemux_8_io_outputs_6_payload_lkIdx[5:0] ), //o
    .io_outputs_6_payload_wLen       (streamDemux_8_io_outputs_6_payload_wLen[2:0]  ), //o
    .io_outputs_7_valid              (streamDemux_8_io_outputs_7_valid              ), //o
    .io_outputs_7_ready              (streamDemux_8_io_outputs_7_ready              ), //i
    .io_outputs_7_payload_nId        (streamDemux_8_io_outputs_7_payload_nId        ), //o
    .io_outputs_7_payload_tId        (streamDemux_8_io_outputs_7_payload_tId[18:0]  ), //o
    .io_outputs_7_payload_tabId      (streamDemux_8_io_outputs_7_payload_tabId[2:0] ), //o
    .io_outputs_7_payload_snId       (streamDemux_8_io_outputs_7_payload_snId       ), //o
    .io_outputs_7_payload_txnId      (streamDemux_8_io_outputs_7_payload_txnId[5:0] ), //o
    .io_outputs_7_payload_lkType     (streamDemux_8_io_outputs_7_payload_lkType[1:0]), //o
    .io_outputs_7_payload_lkRelease  (streamDemux_8_io_outputs_7_payload_lkRelease  ), //o
    .io_outputs_7_payload_txnTimeOut (streamDemux_8_io_outputs_7_payload_txnTimeOut ), //o
    .io_outputs_7_payload_txnAbt     (streamDemux_8_io_outputs_7_payload_txnAbt     ), //o
    .io_outputs_7_payload_lkIdx      (streamDemux_8_io_outputs_7_payload_lkIdx[5:0] ), //o
    .io_outputs_7_payload_wLen       (streamDemux_8_io_outputs_7_payload_wLen[2:0]  )  //o
  );
  StreamArbiter lkRespArb (
    .io_inputs_0_valid             (ltAry_0_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_0_ready             (lkRespArb_io_inputs_0_ready                            ), //o
    .io_inputs_0_payload_nId       (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_0_payload_tId       (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_0_payload_tabId     (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_0_payload_snId      (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_0_payload_txnId     (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_0_payload_lkType    (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_0_payload_lkRelease (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_0_payload_txnAbt    (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_0_payload_lkIdx     (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_0_payload_wLen      (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_0_payload_respType  (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_0_payload_lkWaited  (ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_1_valid             (ltAry_1_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_1_ready             (lkRespArb_io_inputs_1_ready                            ), //o
    .io_inputs_1_payload_nId       (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_1_payload_tId       (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_1_payload_tabId     (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_1_payload_snId      (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_1_payload_txnId     (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_1_payload_lkType    (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_1_payload_lkRelease (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_1_payload_txnAbt    (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_1_payload_lkIdx     (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_1_payload_wLen      (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_1_payload_respType  (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_1_payload_lkWaited  (ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_2_valid             (ltAry_2_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_2_ready             (lkRespArb_io_inputs_2_ready                            ), //o
    .io_inputs_2_payload_nId       (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_2_payload_tId       (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_2_payload_tabId     (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_2_payload_snId      (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_2_payload_txnId     (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_2_payload_lkType    (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_2_payload_lkRelease (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_2_payload_txnAbt    (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_2_payload_lkIdx     (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_2_payload_wLen      (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_2_payload_respType  (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_2_payload_lkWaited  (ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_3_valid             (ltAry_3_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_3_ready             (lkRespArb_io_inputs_3_ready                            ), //o
    .io_inputs_3_payload_nId       (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_3_payload_tId       (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_3_payload_tabId     (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_3_payload_snId      (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_3_payload_txnId     (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_3_payload_lkType    (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_3_payload_lkRelease (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_3_payload_txnAbt    (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_3_payload_lkIdx     (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_3_payload_wLen      (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_3_payload_respType  (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_3_payload_lkWaited  (ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_4_valid             (ltAry_4_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_4_ready             (lkRespArb_io_inputs_4_ready                            ), //o
    .io_inputs_4_payload_nId       (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_4_payload_tId       (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_4_payload_tabId     (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_4_payload_snId      (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_4_payload_txnId     (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_4_payload_lkType    (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_4_payload_lkRelease (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_4_payload_txnAbt    (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_4_payload_lkIdx     (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_4_payload_wLen      (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_4_payload_respType  (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_4_payload_lkWaited  (ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_5_valid             (ltAry_5_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_5_ready             (lkRespArb_io_inputs_5_ready                            ), //o
    .io_inputs_5_payload_nId       (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_5_payload_tId       (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_5_payload_tabId     (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_5_payload_snId      (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_5_payload_txnId     (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_5_payload_lkType    (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_5_payload_lkRelease (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_5_payload_txnAbt    (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_5_payload_lkIdx     (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_5_payload_wLen      (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_5_payload_respType  (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_5_payload_lkWaited  (ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_6_valid             (ltAry_6_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_6_ready             (lkRespArb_io_inputs_6_ready                            ), //o
    .io_inputs_6_payload_nId       (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_6_payload_tId       (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_6_payload_tabId     (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_6_payload_snId      (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_6_payload_txnId     (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_6_payload_lkType    (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_6_payload_lkRelease (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_6_payload_txnAbt    (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_6_payload_lkIdx     (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_6_payload_wLen      (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_6_payload_respType  (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_6_payload_lkWaited  (ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_inputs_7_valid             (ltAry_7_io_lkResp_s2mPipe_m2sPipe_valid                ), //i
    .io_inputs_7_ready             (lkRespArb_io_inputs_7_ready                            ), //o
    .io_inputs_7_payload_nId       (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_nId          ), //i
    .io_inputs_7_payload_tId       (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tId[18:0]    ), //i
    .io_inputs_7_payload_tabId     (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tabId[2:0]   ), //i
    .io_inputs_7_payload_snId      (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_snId         ), //i
    .io_inputs_7_payload_txnId     (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnId[5:0]   ), //i
    .io_inputs_7_payload_lkType    (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType[1:0]  ), //i
    .io_inputs_7_payload_lkRelease (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease    ), //i
    .io_inputs_7_payload_txnAbt    (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt       ), //i
    .io_inputs_7_payload_lkIdx     (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx[5:0]   ), //i
    .io_inputs_7_payload_wLen      (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_wLen[2:0]    ), //i
    .io_inputs_7_payload_respType  (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType[1:0]), //i
    .io_inputs_7_payload_lkWaited  (ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited     ), //i
    .io_output_valid               (lkRespArb_io_output_valid                              ), //o
    .io_output_ready               (lkRespTup_ready                                        ), //i
    .io_output_payload_nId         (lkRespArb_io_output_payload_nId                        ), //o
    .io_output_payload_tId         (lkRespArb_io_output_payload_tId[18:0]                  ), //o
    .io_output_payload_tabId       (lkRespArb_io_output_payload_tabId[2:0]                 ), //o
    .io_output_payload_snId        (lkRespArb_io_output_payload_snId                       ), //o
    .io_output_payload_txnId       (lkRespArb_io_output_payload_txnId[5:0]                 ), //o
    .io_output_payload_lkType      (lkRespArb_io_output_payload_lkType[1:0]                ), //o
    .io_output_payload_lkRelease   (lkRespArb_io_output_payload_lkRelease                  ), //o
    .io_output_payload_txnAbt      (lkRespArb_io_output_payload_txnAbt                     ), //o
    .io_output_payload_lkIdx       (lkRespArb_io_output_payload_lkIdx[5:0]                 ), //o
    .io_output_payload_wLen        (lkRespArb_io_output_payload_wLen[2:0]                  ), //o
    .io_output_payload_respType    (lkRespArb_io_output_payload_respType[1:0]              ), //o
    .io_output_payload_lkWaited    (lkRespArb_io_output_payload_lkWaited                   ), //o
    .io_chosen                     (lkRespArb_io_chosen[2:0]                               ), //o
    .io_chosenOH                   (lkRespArb_io_chosenOH[7:0]                             ), //o
    .clk                           (clk                                                    ), //i
    .resetn                        (resetn                                                 )  //i
  );
  StreamArbiter_1 streamArbiter_8 (
    .io_inputs_0_valid             (lkRespInsTab_valid                             ), //i
    .io_inputs_0_ready             (streamArbiter_8_io_inputs_0_ready              ), //o
    .io_inputs_0_payload_nId       (lkRespInsTab_payload_nId                       ), //i
    .io_inputs_0_payload_tId       (lkRespInsTab_payload_tId[21:0]                 ), //i
    .io_inputs_0_payload_tabId     (lkRespInsTab_payload_tabId[2:0]                ), //i
    .io_inputs_0_payload_snId      (lkRespInsTab_payload_snId                      ), //i
    .io_inputs_0_payload_txnId     (lkRespInsTab_payload_txnId[5:0]                ), //i
    .io_inputs_0_payload_lkType    (lkRespInsTab_payload_lkType[1:0]               ), //i
    .io_inputs_0_payload_lkRelease (lkRespInsTab_payload_lkRelease                 ), //i
    .io_inputs_0_payload_txnAbt    (lkRespInsTab_payload_txnAbt                    ), //i
    .io_inputs_0_payload_lkIdx     (lkRespInsTab_payload_lkIdx[5:0]                ), //i
    .io_inputs_0_payload_wLen      (lkRespInsTab_payload_wLen[2:0]                 ), //i
    .io_inputs_0_payload_respType  (lkRespInsTab_payload_respType[1:0]             ), //i
    .io_inputs_0_payload_lkWaited  (lkRespInsTab_payload_lkWaited                  ), //i
    .io_inputs_1_valid             (lkRespTup_valid                                ), //i
    .io_inputs_1_ready             (streamArbiter_8_io_inputs_1_ready              ), //o
    .io_inputs_1_payload_nId       (lkRespTup_payload_nId                          ), //i
    .io_inputs_1_payload_tId       (lkRespTup_payload_tId[21:0]                    ), //i
    .io_inputs_1_payload_tabId     (lkRespTup_payload_tabId[2:0]                   ), //i
    .io_inputs_1_payload_snId      (lkRespTup_payload_snId                         ), //i
    .io_inputs_1_payload_txnId     (lkRespTup_payload_txnId[5:0]                   ), //i
    .io_inputs_1_payload_lkType    (lkRespTup_payload_lkType[1:0]                  ), //i
    .io_inputs_1_payload_lkRelease (lkRespTup_payload_lkRelease                    ), //i
    .io_inputs_1_payload_txnAbt    (lkRespTup_payload_txnAbt                       ), //i
    .io_inputs_1_payload_lkIdx     (lkRespTup_payload_lkIdx[5:0]                   ), //i
    .io_inputs_1_payload_wLen      (lkRespTup_payload_wLen[2:0]                    ), //i
    .io_inputs_1_payload_respType  (lkRespTup_payload_respType[1:0]                ), //i
    .io_inputs_1_payload_lkWaited  (lkRespTup_payload_lkWaited                     ), //i
    .io_output_valid               (streamArbiter_8_io_output_valid                ), //o
    .io_output_ready               (io_lkResp_ready                                ), //i
    .io_output_payload_nId         (streamArbiter_8_io_output_payload_nId          ), //o
    .io_output_payload_tId         (streamArbiter_8_io_output_payload_tId[21:0]    ), //o
    .io_output_payload_tabId       (streamArbiter_8_io_output_payload_tabId[2:0]   ), //o
    .io_output_payload_snId        (streamArbiter_8_io_output_payload_snId         ), //o
    .io_output_payload_txnId       (streamArbiter_8_io_output_payload_txnId[5:0]   ), //o
    .io_output_payload_lkType      (streamArbiter_8_io_output_payload_lkType[1:0]  ), //o
    .io_output_payload_lkRelease   (streamArbiter_8_io_output_payload_lkRelease    ), //o
    .io_output_payload_txnAbt      (streamArbiter_8_io_output_payload_txnAbt       ), //o
    .io_output_payload_lkIdx       (streamArbiter_8_io_output_payload_lkIdx[5:0]   ), //o
    .io_output_payload_wLen        (streamArbiter_8_io_output_payload_wLen[2:0]    ), //o
    .io_output_payload_respType    (streamArbiter_8_io_output_payload_respType[1:0]), //o
    .io_output_payload_lkWaited    (streamArbiter_8_io_output_payload_lkWaited     ), //o
    .io_chosen                     (streamArbiter_8_io_chosen                      ), //o
    .io_chosenOH                   (streamArbiter_8_io_chosenOH[1:0]               ), //o
    .clk                           (clk                                            ), //i
    .resetn                        (resetn                                         )  //i
  );
  always @(*) begin
    case(streamDemux_7_io_outputs_1_payload_tabId)
      3'b000 : _zz_lkRespInsTab_payload_tId = tupPtr_0;
      3'b001 : _zz_lkRespInsTab_payload_tId = tupPtr_1;
      3'b010 : _zz_lkRespInsTab_payload_tId = tupPtr_2;
      3'b011 : _zz_lkRespInsTab_payload_tId = tupPtr_3;
      3'b100 : _zz_lkRespInsTab_payload_tId = tupPtr_4;
      3'b101 : _zz_lkRespInsTab_payload_tId = tupPtr_5;
      3'b110 : _zz_lkRespInsTab_payload_tId = tupPtr_6;
      default : _zz_lkRespInsTab_payload_tId = tupPtr_7;
    endcase
  end

  always @(*) begin
    case(lkRespInsTab_payload_tabId)
      3'b000 : _zz__zz_tupPtr_0 = tupPtr_0;
      3'b001 : _zz__zz_tupPtr_0 = tupPtr_1;
      3'b010 : _zz__zz_tupPtr_0 = tupPtr_2;
      3'b011 : _zz__zz_tupPtr_0 = tupPtr_3;
      3'b100 : _zz__zz_tupPtr_0 = tupPtr_4;
      3'b101 : _zz__zz_tupPtr_0 = tupPtr_5;
      3'b110 : _zz__zz_tupPtr_0 = tupPtr_6;
      default : _zz__zz_tupPtr_0 = tupPtr_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(lkRespInsTab_payload_lkType)
      LkT_rd : lkRespInsTab_payload_lkType_string = "rd    ";
      LkT_wr : lkRespInsTab_payload_lkType_string = "wr    ";
      LkT_raw : lkRespInsTab_payload_lkType_string = "raw   ";
      LkT_insTab : lkRespInsTab_payload_lkType_string = "insTab";
      default : lkRespInsTab_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkRespInsTab_payload_respType)
      LockRespType_grant : lkRespInsTab_payload_respType_string = "grant    ";
      LockRespType_abort : lkRespInsTab_payload_respType_string = "abort    ";
      LockRespType_waiting : lkRespInsTab_payload_respType_string = "waiting  ";
      LockRespType_release_1 : lkRespInsTab_payload_respType_string = "release_1";
      default : lkRespInsTab_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(lkRespTup_payload_lkType)
      LkT_rd : lkRespTup_payload_lkType_string = "rd    ";
      LkT_wr : lkRespTup_payload_lkType_string = "wr    ";
      LkT_raw : lkRespTup_payload_lkType_string = "raw   ";
      LkT_insTab : lkRespTup_payload_lkType_string = "insTab";
      default : lkRespTup_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(lkRespTup_payload_respType)
      LockRespType_grant : lkRespTup_payload_respType_string = "grant    ";
      LockRespType_abort : lkRespTup_payload_respType_string = "abort    ";
      LockRespType_waiting : lkRespTup_payload_respType_string = "waiting  ";
      LockRespType_release_1 : lkRespTup_payload_respType_string = "release_1";
      default : lkRespTup_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(lkReq2Lt_payload_lkType)
      LkT_rd : lkReq2Lt_payload_lkType_string = "rd    ";
      LkT_wr : lkReq2Lt_payload_lkType_string = "wr    ";
      LkT_raw : lkReq2Lt_payload_lkType_string = "raw   ";
      LkT_insTab : lkReq2Lt_payload_lkType_string = "insTab";
      default : lkReq2Lt_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_0_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_0_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_0_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_0_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_0_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_0_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_0_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_0_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType)
      LkT_rd : _zz_payload_lkType_string = "rd    ";
      LkT_wr : _zz_payload_lkType_string = "wr    ";
      LkT_raw : _zz_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_string = "insTab";
      default : _zz_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_0_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_0_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_1_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_1_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_1_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_1_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_1_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_1_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_1_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_1_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_1)
      LkT_rd : _zz_payload_lkType_1_string = "rd    ";
      LkT_wr : _zz_payload_lkType_1_string = "wr    ";
      LkT_raw : _zz_payload_lkType_1_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_1_string = "insTab";
      default : _zz_payload_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_1_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_1_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_2_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_2_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_2_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_2_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_2_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_2_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_2_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_2_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_2)
      LkT_rd : _zz_payload_lkType_2_string = "rd    ";
      LkT_wr : _zz_payload_lkType_2_string = "wr    ";
      LkT_raw : _zz_payload_lkType_2_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_2_string = "insTab";
      default : _zz_payload_lkType_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_2_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_2_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_3_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_3_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_3_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_3_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_3_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_3_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_3_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_3_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_3)
      LkT_rd : _zz_payload_lkType_3_string = "rd    ";
      LkT_wr : _zz_payload_lkType_3_string = "wr    ";
      LkT_raw : _zz_payload_lkType_3_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_3_string = "insTab";
      default : _zz_payload_lkType_3_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_3_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_3_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_4_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_4_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_4_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_4_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_4_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_4_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_4_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_4_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_4)
      LkT_rd : _zz_payload_lkType_4_string = "rd    ";
      LkT_wr : _zz_payload_lkType_4_string = "wr    ";
      LkT_raw : _zz_payload_lkType_4_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_4_string = "insTab";
      default : _zz_payload_lkType_4_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_4_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_4_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_5_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_5_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_5_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_5_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_5_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_5_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_5_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_5_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_5)
      LkT_rd : _zz_payload_lkType_5_string = "rd    ";
      LkT_wr : _zz_payload_lkType_5_string = "wr    ";
      LkT_raw : _zz_payload_lkType_5_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_5_string = "insTab";
      default : _zz_payload_lkType_5_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_5_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_5_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_6_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_6_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_6_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_6_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_6_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_6_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_6_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_6_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_6)
      LkT_rd : _zz_payload_lkType_6_string = "rd    ";
      LkT_wr : _zz_payload_lkType_6_string = "wr    ";
      LkT_raw : _zz_payload_lkType_6_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_6_string = "insTab";
      default : _zz_payload_lkType_6_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_6_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_6_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_7_s2mPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_7_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_7_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_7_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_7_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_7_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_7_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_7_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_lkType_7)
      LkT_rd : _zz_payload_lkType_7_string = "rd    ";
      LkT_wr : _zz_payload_lkType_7_string = "wr    ";
      LkT_raw : _zz_payload_lkType_7_string = "raw   ";
      LkT_insTab : _zz_payload_lkType_7_string = "insTab";
      default : _zz_payload_lkType_7_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamDemux_8_io_outputs_7_s2mPipe_rData_lkType)
      LkT_rd : streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string = "insTab";
      default : streamDemux_8_io_outputs_7_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_rData_lkType)
      LkT_rd : ltAry_0_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_0_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_0_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_0_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_0_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_0_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_0_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_0_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_0_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_0_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_0_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_0_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_0_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_0_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_0_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_0_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_0_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_0_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_0_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_0_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_0_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_0_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_rData_lkType)
      LkT_rd : ltAry_1_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_1_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_1_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_1_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_1_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_1_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_1_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_1_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_1_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_1_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_1_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_1_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_1_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_1_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_1_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_1_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_1_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_1_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_1_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_1_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_1_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_1_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_rData_lkType)
      LkT_rd : ltAry_2_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_2_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_2_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_2_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_2_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_2_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_2_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_2_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_2_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_2_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_2_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_2_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_2_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_2_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_2_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_2_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_2_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_2_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_2_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_2_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_2_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_2_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_rData_lkType)
      LkT_rd : ltAry_3_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_3_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_3_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_3_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_3_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_3_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_3_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_3_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_3_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_3_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_3_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_3_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_3_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_3_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_3_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_3_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_3_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_3_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_3_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_3_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_3_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_3_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_rData_lkType)
      LkT_rd : ltAry_4_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_4_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_4_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_4_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_4_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_4_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_4_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_4_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_4_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_4_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_4_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_4_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_4_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_4_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_4_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_4_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_4_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_4_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_4_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_4_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_4_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_4_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_rData_lkType)
      LkT_rd : ltAry_5_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_5_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_5_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_5_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_5_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_5_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_5_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_5_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_5_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_5_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_5_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_5_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_5_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_5_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_5_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_5_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_5_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_5_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_5_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_5_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_5_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_5_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_rData_lkType)
      LkT_rd : ltAry_6_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_6_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_6_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_6_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_6_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_6_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_6_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_6_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_6_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_6_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_6_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_6_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_6_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_6_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_6_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_6_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_6_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_6_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_6_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_6_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_6_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_6_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_rData_lkType)
      LkT_rd : ltAry_7_io_lkResp_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_7_io_lkResp_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_7_io_lkResp_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_7_io_lkResp_rData_lkType_string = "insTab";
      default : ltAry_7_io_lkResp_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_rData_respType)
      LockRespType_grant : ltAry_7_io_lkResp_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_7_io_lkResp_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_7_io_lkResp_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_7_io_lkResp_rData_respType_string = "release_1";
      default : ltAry_7_io_lkResp_rData_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType)
      LkT_rd : _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "rd    ";
      LkT_wr : _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "wr    ";
      LkT_raw : _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "insTab";
      default : _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_ltAry_7_io_lkResp_s2mPipe_payload_respType)
      LockRespType_grant : _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "release_1";
      default : _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType)
      LkT_rd : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "rd    ";
      LkT_wr : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "wr    ";
      LkT_raw : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "raw   ";
      LkT_insTab : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "insTab";
      default : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType)
      LockRespType_grant : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "grant    ";
      LockRespType_abort : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "abort    ";
      LockRespType_waiting : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "release_1";
      default : ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_rData_lkType)
      LkT_rd : ltAry_7_io_lkResp_s2mPipe_rData_lkType_string = "rd    ";
      LkT_wr : ltAry_7_io_lkResp_s2mPipe_rData_lkType_string = "wr    ";
      LkT_raw : ltAry_7_io_lkResp_s2mPipe_rData_lkType_string = "raw   ";
      LkT_insTab : ltAry_7_io_lkResp_s2mPipe_rData_lkType_string = "insTab";
      default : ltAry_7_io_lkResp_s2mPipe_rData_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(ltAry_7_io_lkResp_s2mPipe_rData_respType)
      LockRespType_grant : ltAry_7_io_lkResp_s2mPipe_rData_respType_string = "grant    ";
      LockRespType_abort : ltAry_7_io_lkResp_s2mPipe_rData_respType_string = "abort    ";
      LockRespType_waiting : ltAry_7_io_lkResp_s2mPipe_rData_respType_string = "waiting  ";
      LockRespType_release_1 : ltAry_7_io_lkResp_s2mPipe_rData_respType_string = "release_1";
      default : ltAry_7_io_lkResp_s2mPipe_rData_respType_string = "?????????";
    endcase
  end
  `endif

  assign io_lkReq_ready = streamDemux_7_io_input_ready;
  assign streamDemux_7_io_select = ((io_lkReq_payload_lkType == LkT_insTab) ? 1'b1 : 1'b0);
  assign lkRespInsTab_valid = streamDemux_7_io_outputs_1_valid;
  assign lkRespInsTab_payload_nId = streamDemux_7_io_outputs_1_payload_nId;
  always @(*) begin
    lkRespInsTab_payload_tId = streamDemux_7_io_outputs_1_payload_tId;
    lkRespInsTab_payload_tId = _zz_lkRespInsTab_payload_tId;
  end

  assign lkRespInsTab_payload_tabId = streamDemux_7_io_outputs_1_payload_tabId;
  assign lkRespInsTab_payload_snId = streamDemux_7_io_outputs_1_payload_snId;
  assign lkRespInsTab_payload_txnId = streamDemux_7_io_outputs_1_payload_txnId;
  assign lkRespInsTab_payload_lkType = streamDemux_7_io_outputs_1_payload_lkType;
  assign lkRespInsTab_payload_lkRelease = streamDemux_7_io_outputs_1_payload_lkRelease;
  assign lkRespInsTab_payload_txnAbt = streamDemux_7_io_outputs_1_payload_txnAbt;
  assign lkRespInsTab_payload_lkIdx = streamDemux_7_io_outputs_1_payload_lkIdx;
  assign lkRespInsTab_payload_wLen = streamDemux_7_io_outputs_1_payload_wLen;
  assign lkRespInsTab_payload_respType = LockRespType_grant;
  assign lkRespInsTab_payload_lkWaited = 1'b0;
  assign lkRespInsTab_fire = (lkRespInsTab_valid && lkRespInsTab_ready);
  assign _zz_1 = ({7'd0,1'b1} <<< lkRespInsTab_payload_tabId);
  assign _zz_tupPtr_0 = (_zz__zz_tupPtr_0 + streamDemux_7_io_outputs_1_payload_tId);
  assign lkReq2Lt_valid = streamDemux_7_io_outputs_0_valid;
  assign lkReq2Lt_payload_nId = io_lkReq_payload_nId;
  assign lkReq2Lt_payload_tabId = io_lkReq_payload_tabId;
  assign lkReq2Lt_payload_snId = io_lkReq_payload_snId;
  assign lkReq2Lt_payload_txnId = io_lkReq_payload_txnId;
  assign lkReq2Lt_payload_lkType = io_lkReq_payload_lkType;
  assign lkReq2Lt_payload_lkRelease = io_lkReq_payload_lkRelease;
  assign lkReq2Lt_payload_txnTimeOut = io_lkReq_payload_txnTimeOut;
  assign lkReq2Lt_payload_txnAbt = io_lkReq_payload_txnAbt;
  assign lkReq2Lt_payload_lkIdx = io_lkReq_payload_lkIdx;
  assign lkReq2Lt_payload_wLen = io_lkReq_payload_wLen;
  assign lkReq2Lt_payload_tId = {3'd0, _zz_lkReq2Lt_payload_tId};
  assign lkReq2Lt_ready = streamDemux_8_io_input_ready;
  assign streamDemux_8_io_select = io_lkReq_payload_tId[2 : 0];
  assign streamDemux_8_io_outputs_0_ready = (! streamDemux_8_io_outputs_0_rValid);
  assign streamDemux_8_io_outputs_0_s2mPipe_valid = (streamDemux_8_io_outputs_0_valid || streamDemux_8_io_outputs_0_rValid);
  assign _zz_payload_lkType = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_lkType : streamDemux_8_io_outputs_0_payload_lkType);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_nId = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_nId : streamDemux_8_io_outputs_0_payload_nId);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_tId = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_tId : streamDemux_8_io_outputs_0_payload_tId);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_tabId : streamDemux_8_io_outputs_0_payload_tabId);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_snId = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_snId : streamDemux_8_io_outputs_0_payload_snId);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_txnId : streamDemux_8_io_outputs_0_payload_txnId);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_lkType = _zz_payload_lkType;
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_lkRelease : streamDemux_8_io_outputs_0_payload_lkRelease);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_txnTimeOut : streamDemux_8_io_outputs_0_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_txnAbt : streamDemux_8_io_outputs_0_payload_txnAbt);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_lkIdx : streamDemux_8_io_outputs_0_payload_lkIdx);
  assign streamDemux_8_io_outputs_0_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_0_rValid ? streamDemux_8_io_outputs_0_rData_wLen : streamDemux_8_io_outputs_0_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_0_s2mPipe_ready = streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      streamDemux_8_io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_0_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_0_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_0_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_0_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_0_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_0_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_0_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_0_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_0_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_0_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_0_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_0_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_0_s2mPipe_m2sPipe_ready = ltAry_0_io_lkReq_ready;
  assign streamDemux_8_io_outputs_1_ready = (! streamDemux_8_io_outputs_1_rValid);
  assign streamDemux_8_io_outputs_1_s2mPipe_valid = (streamDemux_8_io_outputs_1_valid || streamDemux_8_io_outputs_1_rValid);
  assign _zz_payload_lkType_1 = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_lkType : streamDemux_8_io_outputs_1_payload_lkType);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_nId = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_nId : streamDemux_8_io_outputs_1_payload_nId);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_tId = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_tId : streamDemux_8_io_outputs_1_payload_tId);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_tabId : streamDemux_8_io_outputs_1_payload_tabId);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_snId = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_snId : streamDemux_8_io_outputs_1_payload_snId);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_txnId : streamDemux_8_io_outputs_1_payload_txnId);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_lkType = _zz_payload_lkType_1;
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_lkRelease : streamDemux_8_io_outputs_1_payload_lkRelease);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_txnTimeOut : streamDemux_8_io_outputs_1_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_txnAbt : streamDemux_8_io_outputs_1_payload_txnAbt);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_lkIdx : streamDemux_8_io_outputs_1_payload_lkIdx);
  assign streamDemux_8_io_outputs_1_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_1_rValid ? streamDemux_8_io_outputs_1_rData_wLen : streamDemux_8_io_outputs_1_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_1_s2mPipe_ready = streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_1) begin
      streamDemux_8_io_outputs_1_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_1 = (! streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_1_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_1_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_1_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_1_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_1_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_1_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_1_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_1_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_1_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_1_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_1_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_1_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_1_s2mPipe_m2sPipe_ready = ltAry_1_io_lkReq_ready;
  assign streamDemux_8_io_outputs_2_ready = (! streamDemux_8_io_outputs_2_rValid);
  assign streamDemux_8_io_outputs_2_s2mPipe_valid = (streamDemux_8_io_outputs_2_valid || streamDemux_8_io_outputs_2_rValid);
  assign _zz_payload_lkType_2 = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_lkType : streamDemux_8_io_outputs_2_payload_lkType);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_nId = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_nId : streamDemux_8_io_outputs_2_payload_nId);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_tId = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_tId : streamDemux_8_io_outputs_2_payload_tId);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_tabId : streamDemux_8_io_outputs_2_payload_tabId);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_snId = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_snId : streamDemux_8_io_outputs_2_payload_snId);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_txnId : streamDemux_8_io_outputs_2_payload_txnId);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_lkType = _zz_payload_lkType_2;
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_lkRelease : streamDemux_8_io_outputs_2_payload_lkRelease);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_txnTimeOut : streamDemux_8_io_outputs_2_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_txnAbt : streamDemux_8_io_outputs_2_payload_txnAbt);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_lkIdx : streamDemux_8_io_outputs_2_payload_lkIdx);
  assign streamDemux_8_io_outputs_2_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_2_rValid ? streamDemux_8_io_outputs_2_rData_wLen : streamDemux_8_io_outputs_2_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_2_s2mPipe_ready = streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_2) begin
      streamDemux_8_io_outputs_2_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_2 = (! streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_2_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_2_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_2_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_2_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_2_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_2_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_2_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_2_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_2_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_2_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_2_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_2_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_2_s2mPipe_m2sPipe_ready = ltAry_2_io_lkReq_ready;
  assign streamDemux_8_io_outputs_3_ready = (! streamDemux_8_io_outputs_3_rValid);
  assign streamDemux_8_io_outputs_3_s2mPipe_valid = (streamDemux_8_io_outputs_3_valid || streamDemux_8_io_outputs_3_rValid);
  assign _zz_payload_lkType_3 = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_lkType : streamDemux_8_io_outputs_3_payload_lkType);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_nId = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_nId : streamDemux_8_io_outputs_3_payload_nId);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_tId = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_tId : streamDemux_8_io_outputs_3_payload_tId);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_tabId : streamDemux_8_io_outputs_3_payload_tabId);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_snId = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_snId : streamDemux_8_io_outputs_3_payload_snId);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_txnId : streamDemux_8_io_outputs_3_payload_txnId);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_lkType = _zz_payload_lkType_3;
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_lkRelease : streamDemux_8_io_outputs_3_payload_lkRelease);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_txnTimeOut : streamDemux_8_io_outputs_3_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_txnAbt : streamDemux_8_io_outputs_3_payload_txnAbt);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_lkIdx : streamDemux_8_io_outputs_3_payload_lkIdx);
  assign streamDemux_8_io_outputs_3_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_3_rValid ? streamDemux_8_io_outputs_3_rData_wLen : streamDemux_8_io_outputs_3_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_3_s2mPipe_ready = streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_3) begin
      streamDemux_8_io_outputs_3_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_3 = (! streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_3_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_3_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_3_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_3_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_3_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_3_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_3_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_3_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_3_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_3_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_3_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_3_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_3_s2mPipe_m2sPipe_ready = ltAry_3_io_lkReq_ready;
  assign streamDemux_8_io_outputs_4_ready = (! streamDemux_8_io_outputs_4_rValid);
  assign streamDemux_8_io_outputs_4_s2mPipe_valid = (streamDemux_8_io_outputs_4_valid || streamDemux_8_io_outputs_4_rValid);
  assign _zz_payload_lkType_4 = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_lkType : streamDemux_8_io_outputs_4_payload_lkType);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_nId = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_nId : streamDemux_8_io_outputs_4_payload_nId);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_tId = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_tId : streamDemux_8_io_outputs_4_payload_tId);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_tabId : streamDemux_8_io_outputs_4_payload_tabId);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_snId = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_snId : streamDemux_8_io_outputs_4_payload_snId);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_txnId : streamDemux_8_io_outputs_4_payload_txnId);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_lkType = _zz_payload_lkType_4;
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_lkRelease : streamDemux_8_io_outputs_4_payload_lkRelease);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_txnTimeOut : streamDemux_8_io_outputs_4_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_txnAbt : streamDemux_8_io_outputs_4_payload_txnAbt);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_lkIdx : streamDemux_8_io_outputs_4_payload_lkIdx);
  assign streamDemux_8_io_outputs_4_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_4_rValid ? streamDemux_8_io_outputs_4_rData_wLen : streamDemux_8_io_outputs_4_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_4_s2mPipe_ready = streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_4) begin
      streamDemux_8_io_outputs_4_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_4 = (! streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_4_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_4_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_4_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_4_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_4_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_4_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_4_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_4_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_4_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_4_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_4_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_4_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_4_s2mPipe_m2sPipe_ready = ltAry_4_io_lkReq_ready;
  assign streamDemux_8_io_outputs_5_ready = (! streamDemux_8_io_outputs_5_rValid);
  assign streamDemux_8_io_outputs_5_s2mPipe_valid = (streamDemux_8_io_outputs_5_valid || streamDemux_8_io_outputs_5_rValid);
  assign _zz_payload_lkType_5 = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_lkType : streamDemux_8_io_outputs_5_payload_lkType);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_nId = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_nId : streamDemux_8_io_outputs_5_payload_nId);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_tId = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_tId : streamDemux_8_io_outputs_5_payload_tId);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_tabId : streamDemux_8_io_outputs_5_payload_tabId);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_snId = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_snId : streamDemux_8_io_outputs_5_payload_snId);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_txnId : streamDemux_8_io_outputs_5_payload_txnId);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_lkType = _zz_payload_lkType_5;
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_lkRelease : streamDemux_8_io_outputs_5_payload_lkRelease);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_txnTimeOut : streamDemux_8_io_outputs_5_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_txnAbt : streamDemux_8_io_outputs_5_payload_txnAbt);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_lkIdx : streamDemux_8_io_outputs_5_payload_lkIdx);
  assign streamDemux_8_io_outputs_5_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_5_rValid ? streamDemux_8_io_outputs_5_rData_wLen : streamDemux_8_io_outputs_5_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_5_s2mPipe_ready = streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_5) begin
      streamDemux_8_io_outputs_5_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_5 = (! streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_5_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_5_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_5_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_5_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_5_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_5_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_5_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_5_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_5_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_5_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_5_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_5_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_5_s2mPipe_m2sPipe_ready = ltAry_5_io_lkReq_ready;
  assign streamDemux_8_io_outputs_6_ready = (! streamDemux_8_io_outputs_6_rValid);
  assign streamDemux_8_io_outputs_6_s2mPipe_valid = (streamDemux_8_io_outputs_6_valid || streamDemux_8_io_outputs_6_rValid);
  assign _zz_payload_lkType_6 = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_lkType : streamDemux_8_io_outputs_6_payload_lkType);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_nId = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_nId : streamDemux_8_io_outputs_6_payload_nId);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_tId = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_tId : streamDemux_8_io_outputs_6_payload_tId);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_tabId : streamDemux_8_io_outputs_6_payload_tabId);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_snId = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_snId : streamDemux_8_io_outputs_6_payload_snId);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_txnId : streamDemux_8_io_outputs_6_payload_txnId);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_lkType = _zz_payload_lkType_6;
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_lkRelease : streamDemux_8_io_outputs_6_payload_lkRelease);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_txnTimeOut : streamDemux_8_io_outputs_6_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_txnAbt : streamDemux_8_io_outputs_6_payload_txnAbt);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_lkIdx : streamDemux_8_io_outputs_6_payload_lkIdx);
  assign streamDemux_8_io_outputs_6_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_6_rValid ? streamDemux_8_io_outputs_6_rData_wLen : streamDemux_8_io_outputs_6_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_6_s2mPipe_ready = streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_6) begin
      streamDemux_8_io_outputs_6_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_6 = (! streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_6_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_6_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_6_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_6_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_6_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_6_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_6_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_6_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_6_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_6_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_6_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_6_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_6_s2mPipe_m2sPipe_ready = ltAry_6_io_lkReq_ready;
  assign streamDemux_8_io_outputs_7_ready = (! streamDemux_8_io_outputs_7_rValid);
  assign streamDemux_8_io_outputs_7_s2mPipe_valid = (streamDemux_8_io_outputs_7_valid || streamDemux_8_io_outputs_7_rValid);
  assign _zz_payload_lkType_7 = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_lkType : streamDemux_8_io_outputs_7_payload_lkType);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_nId = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_nId : streamDemux_8_io_outputs_7_payload_nId);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_tId = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_tId : streamDemux_8_io_outputs_7_payload_tId);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_tabId = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_tabId : streamDemux_8_io_outputs_7_payload_tabId);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_snId = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_snId : streamDemux_8_io_outputs_7_payload_snId);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_txnId = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_txnId : streamDemux_8_io_outputs_7_payload_txnId);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_lkType = _zz_payload_lkType_7;
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_lkRelease = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_lkRelease : streamDemux_8_io_outputs_7_payload_lkRelease);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_txnTimeOut = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_txnTimeOut : streamDemux_8_io_outputs_7_payload_txnTimeOut);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_txnAbt = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_txnAbt : streamDemux_8_io_outputs_7_payload_txnAbt);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_lkIdx = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_lkIdx : streamDemux_8_io_outputs_7_payload_lkIdx);
  assign streamDemux_8_io_outputs_7_s2mPipe_payload_wLen = (streamDemux_8_io_outputs_7_rValid ? streamDemux_8_io_outputs_7_rData_wLen : streamDemux_8_io_outputs_7_payload_wLen);
  always @(*) begin
    streamDemux_8_io_outputs_7_s2mPipe_ready = streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_7) begin
      streamDemux_8_io_outputs_7_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_7 = (! streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_valid);
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_valid = streamDemux_8_io_outputs_7_s2mPipe_rValid;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_nId = streamDemux_8_io_outputs_7_s2mPipe_rData_nId;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tId = streamDemux_8_io_outputs_7_s2mPipe_rData_tId;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_tabId = streamDemux_8_io_outputs_7_s2mPipe_rData_tabId;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_snId = streamDemux_8_io_outputs_7_s2mPipe_rData_snId;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnId = streamDemux_8_io_outputs_7_s2mPipe_rData_txnId;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkType = streamDemux_8_io_outputs_7_s2mPipe_rData_lkType;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkRelease = streamDemux_8_io_outputs_7_s2mPipe_rData_lkRelease;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnTimeOut = streamDemux_8_io_outputs_7_s2mPipe_rData_txnTimeOut;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_txnAbt = streamDemux_8_io_outputs_7_s2mPipe_rData_txnAbt;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_lkIdx = streamDemux_8_io_outputs_7_s2mPipe_rData_lkIdx;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_payload_wLen = streamDemux_8_io_outputs_7_s2mPipe_rData_wLen;
  assign streamDemux_8_io_outputs_7_s2mPipe_m2sPipe_ready = ltAry_7_io_lkReq_ready;
  assign ltAry_0_io_lkResp_ready = (! ltAry_0_io_lkResp_rValid);
  assign ltAry_0_io_lkResp_s2mPipe_valid = (ltAry_0_io_lkResp_valid || ltAry_0_io_lkResp_rValid);
  assign _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_lkType : ltAry_0_io_lkResp_payload_lkType);
  assign _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_respType : ltAry_0_io_lkResp_payload_respType);
  assign ltAry_0_io_lkResp_s2mPipe_payload_nId = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_nId : ltAry_0_io_lkResp_payload_nId);
  assign ltAry_0_io_lkResp_s2mPipe_payload_tId = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_tId : ltAry_0_io_lkResp_payload_tId);
  assign ltAry_0_io_lkResp_s2mPipe_payload_tabId = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_tabId : ltAry_0_io_lkResp_payload_tabId);
  assign ltAry_0_io_lkResp_s2mPipe_payload_snId = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_snId : ltAry_0_io_lkResp_payload_snId);
  assign ltAry_0_io_lkResp_s2mPipe_payload_txnId = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_txnId : ltAry_0_io_lkResp_payload_txnId);
  assign ltAry_0_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_0_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_0_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_lkRelease : ltAry_0_io_lkResp_payload_lkRelease);
  assign ltAry_0_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_txnAbt : ltAry_0_io_lkResp_payload_txnAbt);
  assign ltAry_0_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_lkIdx : ltAry_0_io_lkResp_payload_lkIdx);
  assign ltAry_0_io_lkResp_s2mPipe_payload_wLen = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_wLen : ltAry_0_io_lkResp_payload_wLen);
  assign ltAry_0_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_0_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_0_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_0_io_lkResp_rValid ? ltAry_0_io_lkResp_rData_lkWaited : ltAry_0_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_0_io_lkResp_s2mPipe_ready = ltAry_0_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_8) begin
      ltAry_0_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_8 = (! ltAry_0_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_0_io_lkResp_s2mPipe_rValid;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_0_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_0_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_0_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_0_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_0_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_0_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_0_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_0_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_0_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_0_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_0_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_0_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_0_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_0_ready;
  assign ltAry_1_io_lkResp_ready = (! ltAry_1_io_lkResp_rValid);
  assign ltAry_1_io_lkResp_s2mPipe_valid = (ltAry_1_io_lkResp_valid || ltAry_1_io_lkResp_rValid);
  assign _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_lkType : ltAry_1_io_lkResp_payload_lkType);
  assign _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_respType : ltAry_1_io_lkResp_payload_respType);
  assign ltAry_1_io_lkResp_s2mPipe_payload_nId = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_nId : ltAry_1_io_lkResp_payload_nId);
  assign ltAry_1_io_lkResp_s2mPipe_payload_tId = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_tId : ltAry_1_io_lkResp_payload_tId);
  assign ltAry_1_io_lkResp_s2mPipe_payload_tabId = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_tabId : ltAry_1_io_lkResp_payload_tabId);
  assign ltAry_1_io_lkResp_s2mPipe_payload_snId = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_snId : ltAry_1_io_lkResp_payload_snId);
  assign ltAry_1_io_lkResp_s2mPipe_payload_txnId = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_txnId : ltAry_1_io_lkResp_payload_txnId);
  assign ltAry_1_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_1_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_1_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_lkRelease : ltAry_1_io_lkResp_payload_lkRelease);
  assign ltAry_1_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_txnAbt : ltAry_1_io_lkResp_payload_txnAbt);
  assign ltAry_1_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_lkIdx : ltAry_1_io_lkResp_payload_lkIdx);
  assign ltAry_1_io_lkResp_s2mPipe_payload_wLen = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_wLen : ltAry_1_io_lkResp_payload_wLen);
  assign ltAry_1_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_1_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_1_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_1_io_lkResp_rValid ? ltAry_1_io_lkResp_rData_lkWaited : ltAry_1_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_1_io_lkResp_s2mPipe_ready = ltAry_1_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_9) begin
      ltAry_1_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_9 = (! ltAry_1_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_1_io_lkResp_s2mPipe_rValid;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_1_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_1_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_1_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_1_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_1_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_1_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_1_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_1_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_1_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_1_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_1_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_1_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_1_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_1_ready;
  assign ltAry_2_io_lkResp_ready = (! ltAry_2_io_lkResp_rValid);
  assign ltAry_2_io_lkResp_s2mPipe_valid = (ltAry_2_io_lkResp_valid || ltAry_2_io_lkResp_rValid);
  assign _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_lkType : ltAry_2_io_lkResp_payload_lkType);
  assign _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_respType : ltAry_2_io_lkResp_payload_respType);
  assign ltAry_2_io_lkResp_s2mPipe_payload_nId = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_nId : ltAry_2_io_lkResp_payload_nId);
  assign ltAry_2_io_lkResp_s2mPipe_payload_tId = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_tId : ltAry_2_io_lkResp_payload_tId);
  assign ltAry_2_io_lkResp_s2mPipe_payload_tabId = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_tabId : ltAry_2_io_lkResp_payload_tabId);
  assign ltAry_2_io_lkResp_s2mPipe_payload_snId = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_snId : ltAry_2_io_lkResp_payload_snId);
  assign ltAry_2_io_lkResp_s2mPipe_payload_txnId = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_txnId : ltAry_2_io_lkResp_payload_txnId);
  assign ltAry_2_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_2_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_2_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_lkRelease : ltAry_2_io_lkResp_payload_lkRelease);
  assign ltAry_2_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_txnAbt : ltAry_2_io_lkResp_payload_txnAbt);
  assign ltAry_2_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_lkIdx : ltAry_2_io_lkResp_payload_lkIdx);
  assign ltAry_2_io_lkResp_s2mPipe_payload_wLen = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_wLen : ltAry_2_io_lkResp_payload_wLen);
  assign ltAry_2_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_2_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_2_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_2_io_lkResp_rValid ? ltAry_2_io_lkResp_rData_lkWaited : ltAry_2_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_2_io_lkResp_s2mPipe_ready = ltAry_2_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_10) begin
      ltAry_2_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_10 = (! ltAry_2_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_2_io_lkResp_s2mPipe_rValid;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_2_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_2_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_2_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_2_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_2_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_2_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_2_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_2_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_2_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_2_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_2_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_2_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_2_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_2_ready;
  assign ltAry_3_io_lkResp_ready = (! ltAry_3_io_lkResp_rValid);
  assign ltAry_3_io_lkResp_s2mPipe_valid = (ltAry_3_io_lkResp_valid || ltAry_3_io_lkResp_rValid);
  assign _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_lkType : ltAry_3_io_lkResp_payload_lkType);
  assign _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_respType : ltAry_3_io_lkResp_payload_respType);
  assign ltAry_3_io_lkResp_s2mPipe_payload_nId = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_nId : ltAry_3_io_lkResp_payload_nId);
  assign ltAry_3_io_lkResp_s2mPipe_payload_tId = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_tId : ltAry_3_io_lkResp_payload_tId);
  assign ltAry_3_io_lkResp_s2mPipe_payload_tabId = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_tabId : ltAry_3_io_lkResp_payload_tabId);
  assign ltAry_3_io_lkResp_s2mPipe_payload_snId = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_snId : ltAry_3_io_lkResp_payload_snId);
  assign ltAry_3_io_lkResp_s2mPipe_payload_txnId = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_txnId : ltAry_3_io_lkResp_payload_txnId);
  assign ltAry_3_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_3_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_3_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_lkRelease : ltAry_3_io_lkResp_payload_lkRelease);
  assign ltAry_3_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_txnAbt : ltAry_3_io_lkResp_payload_txnAbt);
  assign ltAry_3_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_lkIdx : ltAry_3_io_lkResp_payload_lkIdx);
  assign ltAry_3_io_lkResp_s2mPipe_payload_wLen = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_wLen : ltAry_3_io_lkResp_payload_wLen);
  assign ltAry_3_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_3_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_3_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_3_io_lkResp_rValid ? ltAry_3_io_lkResp_rData_lkWaited : ltAry_3_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_3_io_lkResp_s2mPipe_ready = ltAry_3_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_11) begin
      ltAry_3_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_11 = (! ltAry_3_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_3_io_lkResp_s2mPipe_rValid;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_3_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_3_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_3_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_3_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_3_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_3_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_3_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_3_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_3_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_3_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_3_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_3_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_3_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_3_ready;
  assign ltAry_4_io_lkResp_ready = (! ltAry_4_io_lkResp_rValid);
  assign ltAry_4_io_lkResp_s2mPipe_valid = (ltAry_4_io_lkResp_valid || ltAry_4_io_lkResp_rValid);
  assign _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_lkType : ltAry_4_io_lkResp_payload_lkType);
  assign _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_respType : ltAry_4_io_lkResp_payload_respType);
  assign ltAry_4_io_lkResp_s2mPipe_payload_nId = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_nId : ltAry_4_io_lkResp_payload_nId);
  assign ltAry_4_io_lkResp_s2mPipe_payload_tId = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_tId : ltAry_4_io_lkResp_payload_tId);
  assign ltAry_4_io_lkResp_s2mPipe_payload_tabId = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_tabId : ltAry_4_io_lkResp_payload_tabId);
  assign ltAry_4_io_lkResp_s2mPipe_payload_snId = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_snId : ltAry_4_io_lkResp_payload_snId);
  assign ltAry_4_io_lkResp_s2mPipe_payload_txnId = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_txnId : ltAry_4_io_lkResp_payload_txnId);
  assign ltAry_4_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_4_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_4_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_lkRelease : ltAry_4_io_lkResp_payload_lkRelease);
  assign ltAry_4_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_txnAbt : ltAry_4_io_lkResp_payload_txnAbt);
  assign ltAry_4_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_lkIdx : ltAry_4_io_lkResp_payload_lkIdx);
  assign ltAry_4_io_lkResp_s2mPipe_payload_wLen = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_wLen : ltAry_4_io_lkResp_payload_wLen);
  assign ltAry_4_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_4_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_4_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_4_io_lkResp_rValid ? ltAry_4_io_lkResp_rData_lkWaited : ltAry_4_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_4_io_lkResp_s2mPipe_ready = ltAry_4_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_12) begin
      ltAry_4_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_12 = (! ltAry_4_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_4_io_lkResp_s2mPipe_rValid;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_4_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_4_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_4_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_4_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_4_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_4_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_4_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_4_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_4_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_4_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_4_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_4_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_4_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_4_ready;
  assign ltAry_5_io_lkResp_ready = (! ltAry_5_io_lkResp_rValid);
  assign ltAry_5_io_lkResp_s2mPipe_valid = (ltAry_5_io_lkResp_valid || ltAry_5_io_lkResp_rValid);
  assign _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_lkType : ltAry_5_io_lkResp_payload_lkType);
  assign _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_respType : ltAry_5_io_lkResp_payload_respType);
  assign ltAry_5_io_lkResp_s2mPipe_payload_nId = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_nId : ltAry_5_io_lkResp_payload_nId);
  assign ltAry_5_io_lkResp_s2mPipe_payload_tId = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_tId : ltAry_5_io_lkResp_payload_tId);
  assign ltAry_5_io_lkResp_s2mPipe_payload_tabId = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_tabId : ltAry_5_io_lkResp_payload_tabId);
  assign ltAry_5_io_lkResp_s2mPipe_payload_snId = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_snId : ltAry_5_io_lkResp_payload_snId);
  assign ltAry_5_io_lkResp_s2mPipe_payload_txnId = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_txnId : ltAry_5_io_lkResp_payload_txnId);
  assign ltAry_5_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_5_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_5_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_lkRelease : ltAry_5_io_lkResp_payload_lkRelease);
  assign ltAry_5_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_txnAbt : ltAry_5_io_lkResp_payload_txnAbt);
  assign ltAry_5_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_lkIdx : ltAry_5_io_lkResp_payload_lkIdx);
  assign ltAry_5_io_lkResp_s2mPipe_payload_wLen = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_wLen : ltAry_5_io_lkResp_payload_wLen);
  assign ltAry_5_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_5_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_5_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_5_io_lkResp_rValid ? ltAry_5_io_lkResp_rData_lkWaited : ltAry_5_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_5_io_lkResp_s2mPipe_ready = ltAry_5_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_13) begin
      ltAry_5_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_13 = (! ltAry_5_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_5_io_lkResp_s2mPipe_rValid;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_5_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_5_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_5_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_5_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_5_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_5_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_5_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_5_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_5_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_5_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_5_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_5_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_5_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_5_ready;
  assign ltAry_6_io_lkResp_ready = (! ltAry_6_io_lkResp_rValid);
  assign ltAry_6_io_lkResp_s2mPipe_valid = (ltAry_6_io_lkResp_valid || ltAry_6_io_lkResp_rValid);
  assign _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_lkType : ltAry_6_io_lkResp_payload_lkType);
  assign _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_respType : ltAry_6_io_lkResp_payload_respType);
  assign ltAry_6_io_lkResp_s2mPipe_payload_nId = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_nId : ltAry_6_io_lkResp_payload_nId);
  assign ltAry_6_io_lkResp_s2mPipe_payload_tId = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_tId : ltAry_6_io_lkResp_payload_tId);
  assign ltAry_6_io_lkResp_s2mPipe_payload_tabId = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_tabId : ltAry_6_io_lkResp_payload_tabId);
  assign ltAry_6_io_lkResp_s2mPipe_payload_snId = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_snId : ltAry_6_io_lkResp_payload_snId);
  assign ltAry_6_io_lkResp_s2mPipe_payload_txnId = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_txnId : ltAry_6_io_lkResp_payload_txnId);
  assign ltAry_6_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_6_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_6_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_lkRelease : ltAry_6_io_lkResp_payload_lkRelease);
  assign ltAry_6_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_txnAbt : ltAry_6_io_lkResp_payload_txnAbt);
  assign ltAry_6_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_lkIdx : ltAry_6_io_lkResp_payload_lkIdx);
  assign ltAry_6_io_lkResp_s2mPipe_payload_wLen = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_wLen : ltAry_6_io_lkResp_payload_wLen);
  assign ltAry_6_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_6_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_6_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_6_io_lkResp_rValid ? ltAry_6_io_lkResp_rData_lkWaited : ltAry_6_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_6_io_lkResp_s2mPipe_ready = ltAry_6_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_14) begin
      ltAry_6_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_14 = (! ltAry_6_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_6_io_lkResp_s2mPipe_rValid;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_6_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_6_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_6_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_6_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_6_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_6_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_6_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_6_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_6_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_6_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_6_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_6_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_6_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_6_ready;
  assign ltAry_7_io_lkResp_ready = (! ltAry_7_io_lkResp_rValid);
  assign ltAry_7_io_lkResp_s2mPipe_valid = (ltAry_7_io_lkResp_valid || ltAry_7_io_lkResp_rValid);
  assign _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_lkType : ltAry_7_io_lkResp_payload_lkType);
  assign _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_respType : ltAry_7_io_lkResp_payload_respType);
  assign ltAry_7_io_lkResp_s2mPipe_payload_nId = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_nId : ltAry_7_io_lkResp_payload_nId);
  assign ltAry_7_io_lkResp_s2mPipe_payload_tId = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_tId : ltAry_7_io_lkResp_payload_tId);
  assign ltAry_7_io_lkResp_s2mPipe_payload_tabId = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_tabId : ltAry_7_io_lkResp_payload_tabId);
  assign ltAry_7_io_lkResp_s2mPipe_payload_snId = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_snId : ltAry_7_io_lkResp_payload_snId);
  assign ltAry_7_io_lkResp_s2mPipe_payload_txnId = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_txnId : ltAry_7_io_lkResp_payload_txnId);
  assign ltAry_7_io_lkResp_s2mPipe_payload_lkType = _zz_ltAry_7_io_lkResp_s2mPipe_payload_lkType;
  assign ltAry_7_io_lkResp_s2mPipe_payload_lkRelease = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_lkRelease : ltAry_7_io_lkResp_payload_lkRelease);
  assign ltAry_7_io_lkResp_s2mPipe_payload_txnAbt = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_txnAbt : ltAry_7_io_lkResp_payload_txnAbt);
  assign ltAry_7_io_lkResp_s2mPipe_payload_lkIdx = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_lkIdx : ltAry_7_io_lkResp_payload_lkIdx);
  assign ltAry_7_io_lkResp_s2mPipe_payload_wLen = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_wLen : ltAry_7_io_lkResp_payload_wLen);
  assign ltAry_7_io_lkResp_s2mPipe_payload_respType = _zz_ltAry_7_io_lkResp_s2mPipe_payload_respType;
  assign ltAry_7_io_lkResp_s2mPipe_payload_lkWaited = (ltAry_7_io_lkResp_rValid ? ltAry_7_io_lkResp_rData_lkWaited : ltAry_7_io_lkResp_payload_lkWaited);
  always @(*) begin
    ltAry_7_io_lkResp_s2mPipe_ready = ltAry_7_io_lkResp_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368_15) begin
      ltAry_7_io_lkResp_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368_15 = (! ltAry_7_io_lkResp_s2mPipe_m2sPipe_valid);
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_valid = ltAry_7_io_lkResp_s2mPipe_rValid;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_nId = ltAry_7_io_lkResp_s2mPipe_rData_nId;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tId = ltAry_7_io_lkResp_s2mPipe_rData_tId;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_tabId = ltAry_7_io_lkResp_s2mPipe_rData_tabId;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_snId = ltAry_7_io_lkResp_s2mPipe_rData_snId;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnId = ltAry_7_io_lkResp_s2mPipe_rData_txnId;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkType = ltAry_7_io_lkResp_s2mPipe_rData_lkType;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkRelease = ltAry_7_io_lkResp_s2mPipe_rData_lkRelease;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_txnAbt = ltAry_7_io_lkResp_s2mPipe_rData_txnAbt;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkIdx = ltAry_7_io_lkResp_s2mPipe_rData_lkIdx;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_wLen = ltAry_7_io_lkResp_s2mPipe_rData_wLen;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_respType = ltAry_7_io_lkResp_s2mPipe_rData_respType;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_payload_lkWaited = ltAry_7_io_lkResp_s2mPipe_rData_lkWaited;
  assign ltAry_7_io_lkResp_s2mPipe_m2sPipe_ready = lkRespArb_io_inputs_7_ready;
  assign lkRespTup_valid = lkRespArb_io_output_valid;
  assign lkRespTup_payload_nId = lkRespArb_io_output_payload_nId;
  assign lkRespTup_payload_tabId = lkRespArb_io_output_payload_tabId;
  assign lkRespTup_payload_snId = lkRespArb_io_output_payload_snId;
  assign lkRespTup_payload_txnId = lkRespArb_io_output_payload_txnId;
  assign lkRespTup_payload_lkType = lkRespArb_io_output_payload_lkType;
  assign lkRespTup_payload_lkRelease = lkRespArb_io_output_payload_lkRelease;
  assign lkRespTup_payload_txnAbt = lkRespArb_io_output_payload_txnAbt;
  assign lkRespTup_payload_lkIdx = lkRespArb_io_output_payload_lkIdx;
  assign lkRespTup_payload_wLen = lkRespArb_io_output_payload_wLen;
  assign lkRespTup_payload_respType = lkRespArb_io_output_payload_respType;
  assign lkRespTup_payload_lkWaited = lkRespArb_io_output_payload_lkWaited;
  assign lkRespTup_payload_tId = {lkRespArb_io_output_payload_tId,lkRespArb_io_chosen};
  assign lkRespInsTab_ready = streamArbiter_8_io_inputs_0_ready;
  assign lkRespTup_ready = streamArbiter_8_io_inputs_1_ready;
  assign io_lkResp_valid = streamArbiter_8_io_output_valid;
  assign io_lkResp_payload_nId = streamArbiter_8_io_output_payload_nId;
  assign io_lkResp_payload_tId = streamArbiter_8_io_output_payload_tId;
  assign io_lkResp_payload_tabId = streamArbiter_8_io_output_payload_tabId;
  assign io_lkResp_payload_snId = streamArbiter_8_io_output_payload_snId;
  assign io_lkResp_payload_txnId = streamArbiter_8_io_output_payload_txnId;
  assign io_lkResp_payload_lkType = streamArbiter_8_io_output_payload_lkType;
  assign io_lkResp_payload_lkRelease = streamArbiter_8_io_output_payload_lkRelease;
  assign io_lkResp_payload_txnAbt = streamArbiter_8_io_output_payload_txnAbt;
  assign io_lkResp_payload_lkIdx = streamArbiter_8_io_output_payload_lkIdx;
  assign io_lkResp_payload_wLen = streamArbiter_8_io_output_payload_wLen;
  assign io_lkResp_payload_respType = streamArbiter_8_io_output_payload_respType;
  assign io_lkResp_payload_lkWaited = streamArbiter_8_io_output_payload_lkWaited;
  always @(posedge clk) begin
    if(!resetn) begin
      tupPtr_0 <= 22'h0;
      tupPtr_1 <= 22'h0;
      tupPtr_2 <= 22'h0;
      tupPtr_3 <= 22'h0;
      tupPtr_4 <= 22'h0;
      tupPtr_5 <= 22'h0;
      tupPtr_6 <= 22'h0;
      tupPtr_7 <= 22'h0;
      streamDemux_8_io_outputs_0_rValid <= 1'b0;
      streamDemux_8_io_outputs_0_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_1_rValid <= 1'b0;
      streamDemux_8_io_outputs_1_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_2_rValid <= 1'b0;
      streamDemux_8_io_outputs_2_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_3_rValid <= 1'b0;
      streamDemux_8_io_outputs_3_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_4_rValid <= 1'b0;
      streamDemux_8_io_outputs_4_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_5_rValid <= 1'b0;
      streamDemux_8_io_outputs_5_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_6_rValid <= 1'b0;
      streamDemux_8_io_outputs_6_s2mPipe_rValid <= 1'b0;
      streamDemux_8_io_outputs_7_rValid <= 1'b0;
      streamDemux_8_io_outputs_7_s2mPipe_rValid <= 1'b0;
      ltAry_0_io_lkResp_rValid <= 1'b0;
      ltAry_0_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_1_io_lkResp_rValid <= 1'b0;
      ltAry_1_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_2_io_lkResp_rValid <= 1'b0;
      ltAry_2_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_3_io_lkResp_rValid <= 1'b0;
      ltAry_3_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_4_io_lkResp_rValid <= 1'b0;
      ltAry_4_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_5_io_lkResp_rValid <= 1'b0;
      ltAry_5_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_6_io_lkResp_rValid <= 1'b0;
      ltAry_6_io_lkResp_s2mPipe_rValid <= 1'b0;
      ltAry_7_io_lkResp_rValid <= 1'b0;
      ltAry_7_io_lkResp_s2mPipe_rValid <= 1'b0;
    end else begin
      if(lkRespInsTab_fire) begin
        if(_zz_1[0]) begin
          tupPtr_0 <= _zz_tupPtr_0;
        end
        if(_zz_1[1]) begin
          tupPtr_1 <= _zz_tupPtr_0;
        end
        if(_zz_1[2]) begin
          tupPtr_2 <= _zz_tupPtr_0;
        end
        if(_zz_1[3]) begin
          tupPtr_3 <= _zz_tupPtr_0;
        end
        if(_zz_1[4]) begin
          tupPtr_4 <= _zz_tupPtr_0;
        end
        if(_zz_1[5]) begin
          tupPtr_5 <= _zz_tupPtr_0;
        end
        if(_zz_1[6]) begin
          tupPtr_6 <= _zz_tupPtr_0;
        end
        if(_zz_1[7]) begin
          tupPtr_7 <= _zz_tupPtr_0;
        end
      end
      if(streamDemux_8_io_outputs_0_valid) begin
        streamDemux_8_io_outputs_0_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_0_s2mPipe_ready) begin
        streamDemux_8_io_outputs_0_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_0_s2mPipe_ready) begin
        streamDemux_8_io_outputs_0_s2mPipe_rValid <= streamDemux_8_io_outputs_0_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_1_valid) begin
        streamDemux_8_io_outputs_1_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_1_s2mPipe_ready) begin
        streamDemux_8_io_outputs_1_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_1_s2mPipe_ready) begin
        streamDemux_8_io_outputs_1_s2mPipe_rValid <= streamDemux_8_io_outputs_1_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_2_valid) begin
        streamDemux_8_io_outputs_2_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_2_s2mPipe_ready) begin
        streamDemux_8_io_outputs_2_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_2_s2mPipe_ready) begin
        streamDemux_8_io_outputs_2_s2mPipe_rValid <= streamDemux_8_io_outputs_2_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_3_valid) begin
        streamDemux_8_io_outputs_3_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_3_s2mPipe_ready) begin
        streamDemux_8_io_outputs_3_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_3_s2mPipe_ready) begin
        streamDemux_8_io_outputs_3_s2mPipe_rValid <= streamDemux_8_io_outputs_3_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_4_valid) begin
        streamDemux_8_io_outputs_4_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_4_s2mPipe_ready) begin
        streamDemux_8_io_outputs_4_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_4_s2mPipe_ready) begin
        streamDemux_8_io_outputs_4_s2mPipe_rValid <= streamDemux_8_io_outputs_4_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_5_valid) begin
        streamDemux_8_io_outputs_5_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_5_s2mPipe_ready) begin
        streamDemux_8_io_outputs_5_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_5_s2mPipe_ready) begin
        streamDemux_8_io_outputs_5_s2mPipe_rValid <= streamDemux_8_io_outputs_5_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_6_valid) begin
        streamDemux_8_io_outputs_6_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_6_s2mPipe_ready) begin
        streamDemux_8_io_outputs_6_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_6_s2mPipe_ready) begin
        streamDemux_8_io_outputs_6_s2mPipe_rValid <= streamDemux_8_io_outputs_6_s2mPipe_valid;
      end
      if(streamDemux_8_io_outputs_7_valid) begin
        streamDemux_8_io_outputs_7_rValid <= 1'b1;
      end
      if(streamDemux_8_io_outputs_7_s2mPipe_ready) begin
        streamDemux_8_io_outputs_7_rValid <= 1'b0;
      end
      if(streamDemux_8_io_outputs_7_s2mPipe_ready) begin
        streamDemux_8_io_outputs_7_s2mPipe_rValid <= streamDemux_8_io_outputs_7_s2mPipe_valid;
      end
      if(ltAry_0_io_lkResp_valid) begin
        ltAry_0_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_0_io_lkResp_s2mPipe_ready) begin
        ltAry_0_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_0_io_lkResp_s2mPipe_ready) begin
        ltAry_0_io_lkResp_s2mPipe_rValid <= ltAry_0_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_1_io_lkResp_valid) begin
        ltAry_1_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_1_io_lkResp_s2mPipe_ready) begin
        ltAry_1_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_1_io_lkResp_s2mPipe_ready) begin
        ltAry_1_io_lkResp_s2mPipe_rValid <= ltAry_1_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_2_io_lkResp_valid) begin
        ltAry_2_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_2_io_lkResp_s2mPipe_ready) begin
        ltAry_2_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_2_io_lkResp_s2mPipe_ready) begin
        ltAry_2_io_lkResp_s2mPipe_rValid <= ltAry_2_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_3_io_lkResp_valid) begin
        ltAry_3_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_3_io_lkResp_s2mPipe_ready) begin
        ltAry_3_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_3_io_lkResp_s2mPipe_ready) begin
        ltAry_3_io_lkResp_s2mPipe_rValid <= ltAry_3_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_4_io_lkResp_valid) begin
        ltAry_4_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_4_io_lkResp_s2mPipe_ready) begin
        ltAry_4_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_4_io_lkResp_s2mPipe_ready) begin
        ltAry_4_io_lkResp_s2mPipe_rValid <= ltAry_4_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_5_io_lkResp_valid) begin
        ltAry_5_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_5_io_lkResp_s2mPipe_ready) begin
        ltAry_5_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_5_io_lkResp_s2mPipe_ready) begin
        ltAry_5_io_lkResp_s2mPipe_rValid <= ltAry_5_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_6_io_lkResp_valid) begin
        ltAry_6_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_6_io_lkResp_s2mPipe_ready) begin
        ltAry_6_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_6_io_lkResp_s2mPipe_ready) begin
        ltAry_6_io_lkResp_s2mPipe_rValid <= ltAry_6_io_lkResp_s2mPipe_valid;
      end
      if(ltAry_7_io_lkResp_valid) begin
        ltAry_7_io_lkResp_rValid <= 1'b1;
      end
      if(ltAry_7_io_lkResp_s2mPipe_ready) begin
        ltAry_7_io_lkResp_rValid <= 1'b0;
      end
      if(ltAry_7_io_lkResp_s2mPipe_ready) begin
        ltAry_7_io_lkResp_s2mPipe_rValid <= ltAry_7_io_lkResp_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(streamDemux_8_io_outputs_0_ready) begin
      streamDemux_8_io_outputs_0_rData_nId <= streamDemux_8_io_outputs_0_payload_nId;
      streamDemux_8_io_outputs_0_rData_tId <= streamDemux_8_io_outputs_0_payload_tId;
      streamDemux_8_io_outputs_0_rData_tabId <= streamDemux_8_io_outputs_0_payload_tabId;
      streamDemux_8_io_outputs_0_rData_snId <= streamDemux_8_io_outputs_0_payload_snId;
      streamDemux_8_io_outputs_0_rData_txnId <= streamDemux_8_io_outputs_0_payload_txnId;
      streamDemux_8_io_outputs_0_rData_lkType <= streamDemux_8_io_outputs_0_payload_lkType;
      streamDemux_8_io_outputs_0_rData_lkRelease <= streamDemux_8_io_outputs_0_payload_lkRelease;
      streamDemux_8_io_outputs_0_rData_txnTimeOut <= streamDemux_8_io_outputs_0_payload_txnTimeOut;
      streamDemux_8_io_outputs_0_rData_txnAbt <= streamDemux_8_io_outputs_0_payload_txnAbt;
      streamDemux_8_io_outputs_0_rData_lkIdx <= streamDemux_8_io_outputs_0_payload_lkIdx;
      streamDemux_8_io_outputs_0_rData_wLen <= streamDemux_8_io_outputs_0_payload_wLen;
    end
    if(streamDemux_8_io_outputs_0_s2mPipe_ready) begin
      streamDemux_8_io_outputs_0_s2mPipe_rData_nId <= streamDemux_8_io_outputs_0_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_0_s2mPipe_rData_tId <= streamDemux_8_io_outputs_0_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_0_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_0_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_0_s2mPipe_rData_snId <= streamDemux_8_io_outputs_0_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_0_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_0_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_0_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_0_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_0_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_0_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_0_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_0_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_0_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_0_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_0_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_0_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_0_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_0_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_1_ready) begin
      streamDemux_8_io_outputs_1_rData_nId <= streamDemux_8_io_outputs_1_payload_nId;
      streamDemux_8_io_outputs_1_rData_tId <= streamDemux_8_io_outputs_1_payload_tId;
      streamDemux_8_io_outputs_1_rData_tabId <= streamDemux_8_io_outputs_1_payload_tabId;
      streamDemux_8_io_outputs_1_rData_snId <= streamDemux_8_io_outputs_1_payload_snId;
      streamDemux_8_io_outputs_1_rData_txnId <= streamDemux_8_io_outputs_1_payload_txnId;
      streamDemux_8_io_outputs_1_rData_lkType <= streamDemux_8_io_outputs_1_payload_lkType;
      streamDemux_8_io_outputs_1_rData_lkRelease <= streamDemux_8_io_outputs_1_payload_lkRelease;
      streamDemux_8_io_outputs_1_rData_txnTimeOut <= streamDemux_8_io_outputs_1_payload_txnTimeOut;
      streamDemux_8_io_outputs_1_rData_txnAbt <= streamDemux_8_io_outputs_1_payload_txnAbt;
      streamDemux_8_io_outputs_1_rData_lkIdx <= streamDemux_8_io_outputs_1_payload_lkIdx;
      streamDemux_8_io_outputs_1_rData_wLen <= streamDemux_8_io_outputs_1_payload_wLen;
    end
    if(streamDemux_8_io_outputs_1_s2mPipe_ready) begin
      streamDemux_8_io_outputs_1_s2mPipe_rData_nId <= streamDemux_8_io_outputs_1_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_1_s2mPipe_rData_tId <= streamDemux_8_io_outputs_1_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_1_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_1_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_1_s2mPipe_rData_snId <= streamDemux_8_io_outputs_1_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_1_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_1_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_1_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_1_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_1_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_1_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_1_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_1_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_1_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_1_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_1_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_1_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_1_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_1_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_2_ready) begin
      streamDemux_8_io_outputs_2_rData_nId <= streamDemux_8_io_outputs_2_payload_nId;
      streamDemux_8_io_outputs_2_rData_tId <= streamDemux_8_io_outputs_2_payload_tId;
      streamDemux_8_io_outputs_2_rData_tabId <= streamDemux_8_io_outputs_2_payload_tabId;
      streamDemux_8_io_outputs_2_rData_snId <= streamDemux_8_io_outputs_2_payload_snId;
      streamDemux_8_io_outputs_2_rData_txnId <= streamDemux_8_io_outputs_2_payload_txnId;
      streamDemux_8_io_outputs_2_rData_lkType <= streamDemux_8_io_outputs_2_payload_lkType;
      streamDemux_8_io_outputs_2_rData_lkRelease <= streamDemux_8_io_outputs_2_payload_lkRelease;
      streamDemux_8_io_outputs_2_rData_txnTimeOut <= streamDemux_8_io_outputs_2_payload_txnTimeOut;
      streamDemux_8_io_outputs_2_rData_txnAbt <= streamDemux_8_io_outputs_2_payload_txnAbt;
      streamDemux_8_io_outputs_2_rData_lkIdx <= streamDemux_8_io_outputs_2_payload_lkIdx;
      streamDemux_8_io_outputs_2_rData_wLen <= streamDemux_8_io_outputs_2_payload_wLen;
    end
    if(streamDemux_8_io_outputs_2_s2mPipe_ready) begin
      streamDemux_8_io_outputs_2_s2mPipe_rData_nId <= streamDemux_8_io_outputs_2_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_2_s2mPipe_rData_tId <= streamDemux_8_io_outputs_2_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_2_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_2_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_2_s2mPipe_rData_snId <= streamDemux_8_io_outputs_2_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_2_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_2_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_2_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_2_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_2_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_2_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_2_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_2_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_2_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_2_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_2_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_2_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_2_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_2_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_3_ready) begin
      streamDemux_8_io_outputs_3_rData_nId <= streamDemux_8_io_outputs_3_payload_nId;
      streamDemux_8_io_outputs_3_rData_tId <= streamDemux_8_io_outputs_3_payload_tId;
      streamDemux_8_io_outputs_3_rData_tabId <= streamDemux_8_io_outputs_3_payload_tabId;
      streamDemux_8_io_outputs_3_rData_snId <= streamDemux_8_io_outputs_3_payload_snId;
      streamDemux_8_io_outputs_3_rData_txnId <= streamDemux_8_io_outputs_3_payload_txnId;
      streamDemux_8_io_outputs_3_rData_lkType <= streamDemux_8_io_outputs_3_payload_lkType;
      streamDemux_8_io_outputs_3_rData_lkRelease <= streamDemux_8_io_outputs_3_payload_lkRelease;
      streamDemux_8_io_outputs_3_rData_txnTimeOut <= streamDemux_8_io_outputs_3_payload_txnTimeOut;
      streamDemux_8_io_outputs_3_rData_txnAbt <= streamDemux_8_io_outputs_3_payload_txnAbt;
      streamDemux_8_io_outputs_3_rData_lkIdx <= streamDemux_8_io_outputs_3_payload_lkIdx;
      streamDemux_8_io_outputs_3_rData_wLen <= streamDemux_8_io_outputs_3_payload_wLen;
    end
    if(streamDemux_8_io_outputs_3_s2mPipe_ready) begin
      streamDemux_8_io_outputs_3_s2mPipe_rData_nId <= streamDemux_8_io_outputs_3_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_3_s2mPipe_rData_tId <= streamDemux_8_io_outputs_3_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_3_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_3_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_3_s2mPipe_rData_snId <= streamDemux_8_io_outputs_3_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_3_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_3_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_3_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_3_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_3_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_3_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_3_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_3_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_3_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_3_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_3_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_3_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_3_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_3_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_4_ready) begin
      streamDemux_8_io_outputs_4_rData_nId <= streamDemux_8_io_outputs_4_payload_nId;
      streamDemux_8_io_outputs_4_rData_tId <= streamDemux_8_io_outputs_4_payload_tId;
      streamDemux_8_io_outputs_4_rData_tabId <= streamDemux_8_io_outputs_4_payload_tabId;
      streamDemux_8_io_outputs_4_rData_snId <= streamDemux_8_io_outputs_4_payload_snId;
      streamDemux_8_io_outputs_4_rData_txnId <= streamDemux_8_io_outputs_4_payload_txnId;
      streamDemux_8_io_outputs_4_rData_lkType <= streamDemux_8_io_outputs_4_payload_lkType;
      streamDemux_8_io_outputs_4_rData_lkRelease <= streamDemux_8_io_outputs_4_payload_lkRelease;
      streamDemux_8_io_outputs_4_rData_txnTimeOut <= streamDemux_8_io_outputs_4_payload_txnTimeOut;
      streamDemux_8_io_outputs_4_rData_txnAbt <= streamDemux_8_io_outputs_4_payload_txnAbt;
      streamDemux_8_io_outputs_4_rData_lkIdx <= streamDemux_8_io_outputs_4_payload_lkIdx;
      streamDemux_8_io_outputs_4_rData_wLen <= streamDemux_8_io_outputs_4_payload_wLen;
    end
    if(streamDemux_8_io_outputs_4_s2mPipe_ready) begin
      streamDemux_8_io_outputs_4_s2mPipe_rData_nId <= streamDemux_8_io_outputs_4_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_4_s2mPipe_rData_tId <= streamDemux_8_io_outputs_4_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_4_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_4_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_4_s2mPipe_rData_snId <= streamDemux_8_io_outputs_4_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_4_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_4_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_4_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_4_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_4_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_4_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_4_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_4_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_4_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_4_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_4_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_4_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_4_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_4_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_5_ready) begin
      streamDemux_8_io_outputs_5_rData_nId <= streamDemux_8_io_outputs_5_payload_nId;
      streamDemux_8_io_outputs_5_rData_tId <= streamDemux_8_io_outputs_5_payload_tId;
      streamDemux_8_io_outputs_5_rData_tabId <= streamDemux_8_io_outputs_5_payload_tabId;
      streamDemux_8_io_outputs_5_rData_snId <= streamDemux_8_io_outputs_5_payload_snId;
      streamDemux_8_io_outputs_5_rData_txnId <= streamDemux_8_io_outputs_5_payload_txnId;
      streamDemux_8_io_outputs_5_rData_lkType <= streamDemux_8_io_outputs_5_payload_lkType;
      streamDemux_8_io_outputs_5_rData_lkRelease <= streamDemux_8_io_outputs_5_payload_lkRelease;
      streamDemux_8_io_outputs_5_rData_txnTimeOut <= streamDemux_8_io_outputs_5_payload_txnTimeOut;
      streamDemux_8_io_outputs_5_rData_txnAbt <= streamDemux_8_io_outputs_5_payload_txnAbt;
      streamDemux_8_io_outputs_5_rData_lkIdx <= streamDemux_8_io_outputs_5_payload_lkIdx;
      streamDemux_8_io_outputs_5_rData_wLen <= streamDemux_8_io_outputs_5_payload_wLen;
    end
    if(streamDemux_8_io_outputs_5_s2mPipe_ready) begin
      streamDemux_8_io_outputs_5_s2mPipe_rData_nId <= streamDemux_8_io_outputs_5_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_5_s2mPipe_rData_tId <= streamDemux_8_io_outputs_5_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_5_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_5_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_5_s2mPipe_rData_snId <= streamDemux_8_io_outputs_5_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_5_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_5_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_5_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_5_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_5_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_5_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_5_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_5_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_5_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_5_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_5_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_5_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_5_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_5_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_6_ready) begin
      streamDemux_8_io_outputs_6_rData_nId <= streamDemux_8_io_outputs_6_payload_nId;
      streamDemux_8_io_outputs_6_rData_tId <= streamDemux_8_io_outputs_6_payload_tId;
      streamDemux_8_io_outputs_6_rData_tabId <= streamDemux_8_io_outputs_6_payload_tabId;
      streamDemux_8_io_outputs_6_rData_snId <= streamDemux_8_io_outputs_6_payload_snId;
      streamDemux_8_io_outputs_6_rData_txnId <= streamDemux_8_io_outputs_6_payload_txnId;
      streamDemux_8_io_outputs_6_rData_lkType <= streamDemux_8_io_outputs_6_payload_lkType;
      streamDemux_8_io_outputs_6_rData_lkRelease <= streamDemux_8_io_outputs_6_payload_lkRelease;
      streamDemux_8_io_outputs_6_rData_txnTimeOut <= streamDemux_8_io_outputs_6_payload_txnTimeOut;
      streamDemux_8_io_outputs_6_rData_txnAbt <= streamDemux_8_io_outputs_6_payload_txnAbt;
      streamDemux_8_io_outputs_6_rData_lkIdx <= streamDemux_8_io_outputs_6_payload_lkIdx;
      streamDemux_8_io_outputs_6_rData_wLen <= streamDemux_8_io_outputs_6_payload_wLen;
    end
    if(streamDemux_8_io_outputs_6_s2mPipe_ready) begin
      streamDemux_8_io_outputs_6_s2mPipe_rData_nId <= streamDemux_8_io_outputs_6_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_6_s2mPipe_rData_tId <= streamDemux_8_io_outputs_6_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_6_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_6_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_6_s2mPipe_rData_snId <= streamDemux_8_io_outputs_6_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_6_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_6_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_6_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_6_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_6_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_6_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_6_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_6_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_6_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_6_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_6_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_6_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_6_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_6_s2mPipe_payload_wLen;
    end
    if(streamDemux_8_io_outputs_7_ready) begin
      streamDemux_8_io_outputs_7_rData_nId <= streamDemux_8_io_outputs_7_payload_nId;
      streamDemux_8_io_outputs_7_rData_tId <= streamDemux_8_io_outputs_7_payload_tId;
      streamDemux_8_io_outputs_7_rData_tabId <= streamDemux_8_io_outputs_7_payload_tabId;
      streamDemux_8_io_outputs_7_rData_snId <= streamDemux_8_io_outputs_7_payload_snId;
      streamDemux_8_io_outputs_7_rData_txnId <= streamDemux_8_io_outputs_7_payload_txnId;
      streamDemux_8_io_outputs_7_rData_lkType <= streamDemux_8_io_outputs_7_payload_lkType;
      streamDemux_8_io_outputs_7_rData_lkRelease <= streamDemux_8_io_outputs_7_payload_lkRelease;
      streamDemux_8_io_outputs_7_rData_txnTimeOut <= streamDemux_8_io_outputs_7_payload_txnTimeOut;
      streamDemux_8_io_outputs_7_rData_txnAbt <= streamDemux_8_io_outputs_7_payload_txnAbt;
      streamDemux_8_io_outputs_7_rData_lkIdx <= streamDemux_8_io_outputs_7_payload_lkIdx;
      streamDemux_8_io_outputs_7_rData_wLen <= streamDemux_8_io_outputs_7_payload_wLen;
    end
    if(streamDemux_8_io_outputs_7_s2mPipe_ready) begin
      streamDemux_8_io_outputs_7_s2mPipe_rData_nId <= streamDemux_8_io_outputs_7_s2mPipe_payload_nId;
      streamDemux_8_io_outputs_7_s2mPipe_rData_tId <= streamDemux_8_io_outputs_7_s2mPipe_payload_tId;
      streamDemux_8_io_outputs_7_s2mPipe_rData_tabId <= streamDemux_8_io_outputs_7_s2mPipe_payload_tabId;
      streamDemux_8_io_outputs_7_s2mPipe_rData_snId <= streamDemux_8_io_outputs_7_s2mPipe_payload_snId;
      streamDemux_8_io_outputs_7_s2mPipe_rData_txnId <= streamDemux_8_io_outputs_7_s2mPipe_payload_txnId;
      streamDemux_8_io_outputs_7_s2mPipe_rData_lkType <= streamDemux_8_io_outputs_7_s2mPipe_payload_lkType;
      streamDemux_8_io_outputs_7_s2mPipe_rData_lkRelease <= streamDemux_8_io_outputs_7_s2mPipe_payload_lkRelease;
      streamDemux_8_io_outputs_7_s2mPipe_rData_txnTimeOut <= streamDemux_8_io_outputs_7_s2mPipe_payload_txnTimeOut;
      streamDemux_8_io_outputs_7_s2mPipe_rData_txnAbt <= streamDemux_8_io_outputs_7_s2mPipe_payload_txnAbt;
      streamDemux_8_io_outputs_7_s2mPipe_rData_lkIdx <= streamDemux_8_io_outputs_7_s2mPipe_payload_lkIdx;
      streamDemux_8_io_outputs_7_s2mPipe_rData_wLen <= streamDemux_8_io_outputs_7_s2mPipe_payload_wLen;
    end
    if(ltAry_0_io_lkResp_ready) begin
      ltAry_0_io_lkResp_rData_nId <= ltAry_0_io_lkResp_payload_nId;
      ltAry_0_io_lkResp_rData_tId <= ltAry_0_io_lkResp_payload_tId;
      ltAry_0_io_lkResp_rData_tabId <= ltAry_0_io_lkResp_payload_tabId;
      ltAry_0_io_lkResp_rData_snId <= ltAry_0_io_lkResp_payload_snId;
      ltAry_0_io_lkResp_rData_txnId <= ltAry_0_io_lkResp_payload_txnId;
      ltAry_0_io_lkResp_rData_lkType <= ltAry_0_io_lkResp_payload_lkType;
      ltAry_0_io_lkResp_rData_lkRelease <= ltAry_0_io_lkResp_payload_lkRelease;
      ltAry_0_io_lkResp_rData_txnAbt <= ltAry_0_io_lkResp_payload_txnAbt;
      ltAry_0_io_lkResp_rData_lkIdx <= ltAry_0_io_lkResp_payload_lkIdx;
      ltAry_0_io_lkResp_rData_wLen <= ltAry_0_io_lkResp_payload_wLen;
      ltAry_0_io_lkResp_rData_respType <= ltAry_0_io_lkResp_payload_respType;
      ltAry_0_io_lkResp_rData_lkWaited <= ltAry_0_io_lkResp_payload_lkWaited;
    end
    if(ltAry_0_io_lkResp_s2mPipe_ready) begin
      ltAry_0_io_lkResp_s2mPipe_rData_nId <= ltAry_0_io_lkResp_s2mPipe_payload_nId;
      ltAry_0_io_lkResp_s2mPipe_rData_tId <= ltAry_0_io_lkResp_s2mPipe_payload_tId;
      ltAry_0_io_lkResp_s2mPipe_rData_tabId <= ltAry_0_io_lkResp_s2mPipe_payload_tabId;
      ltAry_0_io_lkResp_s2mPipe_rData_snId <= ltAry_0_io_lkResp_s2mPipe_payload_snId;
      ltAry_0_io_lkResp_s2mPipe_rData_txnId <= ltAry_0_io_lkResp_s2mPipe_payload_txnId;
      ltAry_0_io_lkResp_s2mPipe_rData_lkType <= ltAry_0_io_lkResp_s2mPipe_payload_lkType;
      ltAry_0_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_0_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_0_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_0_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_0_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_0_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_0_io_lkResp_s2mPipe_rData_wLen <= ltAry_0_io_lkResp_s2mPipe_payload_wLen;
      ltAry_0_io_lkResp_s2mPipe_rData_respType <= ltAry_0_io_lkResp_s2mPipe_payload_respType;
      ltAry_0_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_0_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_1_io_lkResp_ready) begin
      ltAry_1_io_lkResp_rData_nId <= ltAry_1_io_lkResp_payload_nId;
      ltAry_1_io_lkResp_rData_tId <= ltAry_1_io_lkResp_payload_tId;
      ltAry_1_io_lkResp_rData_tabId <= ltAry_1_io_lkResp_payload_tabId;
      ltAry_1_io_lkResp_rData_snId <= ltAry_1_io_lkResp_payload_snId;
      ltAry_1_io_lkResp_rData_txnId <= ltAry_1_io_lkResp_payload_txnId;
      ltAry_1_io_lkResp_rData_lkType <= ltAry_1_io_lkResp_payload_lkType;
      ltAry_1_io_lkResp_rData_lkRelease <= ltAry_1_io_lkResp_payload_lkRelease;
      ltAry_1_io_lkResp_rData_txnAbt <= ltAry_1_io_lkResp_payload_txnAbt;
      ltAry_1_io_lkResp_rData_lkIdx <= ltAry_1_io_lkResp_payload_lkIdx;
      ltAry_1_io_lkResp_rData_wLen <= ltAry_1_io_lkResp_payload_wLen;
      ltAry_1_io_lkResp_rData_respType <= ltAry_1_io_lkResp_payload_respType;
      ltAry_1_io_lkResp_rData_lkWaited <= ltAry_1_io_lkResp_payload_lkWaited;
    end
    if(ltAry_1_io_lkResp_s2mPipe_ready) begin
      ltAry_1_io_lkResp_s2mPipe_rData_nId <= ltAry_1_io_lkResp_s2mPipe_payload_nId;
      ltAry_1_io_lkResp_s2mPipe_rData_tId <= ltAry_1_io_lkResp_s2mPipe_payload_tId;
      ltAry_1_io_lkResp_s2mPipe_rData_tabId <= ltAry_1_io_lkResp_s2mPipe_payload_tabId;
      ltAry_1_io_lkResp_s2mPipe_rData_snId <= ltAry_1_io_lkResp_s2mPipe_payload_snId;
      ltAry_1_io_lkResp_s2mPipe_rData_txnId <= ltAry_1_io_lkResp_s2mPipe_payload_txnId;
      ltAry_1_io_lkResp_s2mPipe_rData_lkType <= ltAry_1_io_lkResp_s2mPipe_payload_lkType;
      ltAry_1_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_1_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_1_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_1_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_1_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_1_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_1_io_lkResp_s2mPipe_rData_wLen <= ltAry_1_io_lkResp_s2mPipe_payload_wLen;
      ltAry_1_io_lkResp_s2mPipe_rData_respType <= ltAry_1_io_lkResp_s2mPipe_payload_respType;
      ltAry_1_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_1_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_2_io_lkResp_ready) begin
      ltAry_2_io_lkResp_rData_nId <= ltAry_2_io_lkResp_payload_nId;
      ltAry_2_io_lkResp_rData_tId <= ltAry_2_io_lkResp_payload_tId;
      ltAry_2_io_lkResp_rData_tabId <= ltAry_2_io_lkResp_payload_tabId;
      ltAry_2_io_lkResp_rData_snId <= ltAry_2_io_lkResp_payload_snId;
      ltAry_2_io_lkResp_rData_txnId <= ltAry_2_io_lkResp_payload_txnId;
      ltAry_2_io_lkResp_rData_lkType <= ltAry_2_io_lkResp_payload_lkType;
      ltAry_2_io_lkResp_rData_lkRelease <= ltAry_2_io_lkResp_payload_lkRelease;
      ltAry_2_io_lkResp_rData_txnAbt <= ltAry_2_io_lkResp_payload_txnAbt;
      ltAry_2_io_lkResp_rData_lkIdx <= ltAry_2_io_lkResp_payload_lkIdx;
      ltAry_2_io_lkResp_rData_wLen <= ltAry_2_io_lkResp_payload_wLen;
      ltAry_2_io_lkResp_rData_respType <= ltAry_2_io_lkResp_payload_respType;
      ltAry_2_io_lkResp_rData_lkWaited <= ltAry_2_io_lkResp_payload_lkWaited;
    end
    if(ltAry_2_io_lkResp_s2mPipe_ready) begin
      ltAry_2_io_lkResp_s2mPipe_rData_nId <= ltAry_2_io_lkResp_s2mPipe_payload_nId;
      ltAry_2_io_lkResp_s2mPipe_rData_tId <= ltAry_2_io_lkResp_s2mPipe_payload_tId;
      ltAry_2_io_lkResp_s2mPipe_rData_tabId <= ltAry_2_io_lkResp_s2mPipe_payload_tabId;
      ltAry_2_io_lkResp_s2mPipe_rData_snId <= ltAry_2_io_lkResp_s2mPipe_payload_snId;
      ltAry_2_io_lkResp_s2mPipe_rData_txnId <= ltAry_2_io_lkResp_s2mPipe_payload_txnId;
      ltAry_2_io_lkResp_s2mPipe_rData_lkType <= ltAry_2_io_lkResp_s2mPipe_payload_lkType;
      ltAry_2_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_2_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_2_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_2_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_2_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_2_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_2_io_lkResp_s2mPipe_rData_wLen <= ltAry_2_io_lkResp_s2mPipe_payload_wLen;
      ltAry_2_io_lkResp_s2mPipe_rData_respType <= ltAry_2_io_lkResp_s2mPipe_payload_respType;
      ltAry_2_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_2_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_3_io_lkResp_ready) begin
      ltAry_3_io_lkResp_rData_nId <= ltAry_3_io_lkResp_payload_nId;
      ltAry_3_io_lkResp_rData_tId <= ltAry_3_io_lkResp_payload_tId;
      ltAry_3_io_lkResp_rData_tabId <= ltAry_3_io_lkResp_payload_tabId;
      ltAry_3_io_lkResp_rData_snId <= ltAry_3_io_lkResp_payload_snId;
      ltAry_3_io_lkResp_rData_txnId <= ltAry_3_io_lkResp_payload_txnId;
      ltAry_3_io_lkResp_rData_lkType <= ltAry_3_io_lkResp_payload_lkType;
      ltAry_3_io_lkResp_rData_lkRelease <= ltAry_3_io_lkResp_payload_lkRelease;
      ltAry_3_io_lkResp_rData_txnAbt <= ltAry_3_io_lkResp_payload_txnAbt;
      ltAry_3_io_lkResp_rData_lkIdx <= ltAry_3_io_lkResp_payload_lkIdx;
      ltAry_3_io_lkResp_rData_wLen <= ltAry_3_io_lkResp_payload_wLen;
      ltAry_3_io_lkResp_rData_respType <= ltAry_3_io_lkResp_payload_respType;
      ltAry_3_io_lkResp_rData_lkWaited <= ltAry_3_io_lkResp_payload_lkWaited;
    end
    if(ltAry_3_io_lkResp_s2mPipe_ready) begin
      ltAry_3_io_lkResp_s2mPipe_rData_nId <= ltAry_3_io_lkResp_s2mPipe_payload_nId;
      ltAry_3_io_lkResp_s2mPipe_rData_tId <= ltAry_3_io_lkResp_s2mPipe_payload_tId;
      ltAry_3_io_lkResp_s2mPipe_rData_tabId <= ltAry_3_io_lkResp_s2mPipe_payload_tabId;
      ltAry_3_io_lkResp_s2mPipe_rData_snId <= ltAry_3_io_lkResp_s2mPipe_payload_snId;
      ltAry_3_io_lkResp_s2mPipe_rData_txnId <= ltAry_3_io_lkResp_s2mPipe_payload_txnId;
      ltAry_3_io_lkResp_s2mPipe_rData_lkType <= ltAry_3_io_lkResp_s2mPipe_payload_lkType;
      ltAry_3_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_3_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_3_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_3_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_3_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_3_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_3_io_lkResp_s2mPipe_rData_wLen <= ltAry_3_io_lkResp_s2mPipe_payload_wLen;
      ltAry_3_io_lkResp_s2mPipe_rData_respType <= ltAry_3_io_lkResp_s2mPipe_payload_respType;
      ltAry_3_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_3_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_4_io_lkResp_ready) begin
      ltAry_4_io_lkResp_rData_nId <= ltAry_4_io_lkResp_payload_nId;
      ltAry_4_io_lkResp_rData_tId <= ltAry_4_io_lkResp_payload_tId;
      ltAry_4_io_lkResp_rData_tabId <= ltAry_4_io_lkResp_payload_tabId;
      ltAry_4_io_lkResp_rData_snId <= ltAry_4_io_lkResp_payload_snId;
      ltAry_4_io_lkResp_rData_txnId <= ltAry_4_io_lkResp_payload_txnId;
      ltAry_4_io_lkResp_rData_lkType <= ltAry_4_io_lkResp_payload_lkType;
      ltAry_4_io_lkResp_rData_lkRelease <= ltAry_4_io_lkResp_payload_lkRelease;
      ltAry_4_io_lkResp_rData_txnAbt <= ltAry_4_io_lkResp_payload_txnAbt;
      ltAry_4_io_lkResp_rData_lkIdx <= ltAry_4_io_lkResp_payload_lkIdx;
      ltAry_4_io_lkResp_rData_wLen <= ltAry_4_io_lkResp_payload_wLen;
      ltAry_4_io_lkResp_rData_respType <= ltAry_4_io_lkResp_payload_respType;
      ltAry_4_io_lkResp_rData_lkWaited <= ltAry_4_io_lkResp_payload_lkWaited;
    end
    if(ltAry_4_io_lkResp_s2mPipe_ready) begin
      ltAry_4_io_lkResp_s2mPipe_rData_nId <= ltAry_4_io_lkResp_s2mPipe_payload_nId;
      ltAry_4_io_lkResp_s2mPipe_rData_tId <= ltAry_4_io_lkResp_s2mPipe_payload_tId;
      ltAry_4_io_lkResp_s2mPipe_rData_tabId <= ltAry_4_io_lkResp_s2mPipe_payload_tabId;
      ltAry_4_io_lkResp_s2mPipe_rData_snId <= ltAry_4_io_lkResp_s2mPipe_payload_snId;
      ltAry_4_io_lkResp_s2mPipe_rData_txnId <= ltAry_4_io_lkResp_s2mPipe_payload_txnId;
      ltAry_4_io_lkResp_s2mPipe_rData_lkType <= ltAry_4_io_lkResp_s2mPipe_payload_lkType;
      ltAry_4_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_4_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_4_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_4_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_4_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_4_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_4_io_lkResp_s2mPipe_rData_wLen <= ltAry_4_io_lkResp_s2mPipe_payload_wLen;
      ltAry_4_io_lkResp_s2mPipe_rData_respType <= ltAry_4_io_lkResp_s2mPipe_payload_respType;
      ltAry_4_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_4_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_5_io_lkResp_ready) begin
      ltAry_5_io_lkResp_rData_nId <= ltAry_5_io_lkResp_payload_nId;
      ltAry_5_io_lkResp_rData_tId <= ltAry_5_io_lkResp_payload_tId;
      ltAry_5_io_lkResp_rData_tabId <= ltAry_5_io_lkResp_payload_tabId;
      ltAry_5_io_lkResp_rData_snId <= ltAry_5_io_lkResp_payload_snId;
      ltAry_5_io_lkResp_rData_txnId <= ltAry_5_io_lkResp_payload_txnId;
      ltAry_5_io_lkResp_rData_lkType <= ltAry_5_io_lkResp_payload_lkType;
      ltAry_5_io_lkResp_rData_lkRelease <= ltAry_5_io_lkResp_payload_lkRelease;
      ltAry_5_io_lkResp_rData_txnAbt <= ltAry_5_io_lkResp_payload_txnAbt;
      ltAry_5_io_lkResp_rData_lkIdx <= ltAry_5_io_lkResp_payload_lkIdx;
      ltAry_5_io_lkResp_rData_wLen <= ltAry_5_io_lkResp_payload_wLen;
      ltAry_5_io_lkResp_rData_respType <= ltAry_5_io_lkResp_payload_respType;
      ltAry_5_io_lkResp_rData_lkWaited <= ltAry_5_io_lkResp_payload_lkWaited;
    end
    if(ltAry_5_io_lkResp_s2mPipe_ready) begin
      ltAry_5_io_lkResp_s2mPipe_rData_nId <= ltAry_5_io_lkResp_s2mPipe_payload_nId;
      ltAry_5_io_lkResp_s2mPipe_rData_tId <= ltAry_5_io_lkResp_s2mPipe_payload_tId;
      ltAry_5_io_lkResp_s2mPipe_rData_tabId <= ltAry_5_io_lkResp_s2mPipe_payload_tabId;
      ltAry_5_io_lkResp_s2mPipe_rData_snId <= ltAry_5_io_lkResp_s2mPipe_payload_snId;
      ltAry_5_io_lkResp_s2mPipe_rData_txnId <= ltAry_5_io_lkResp_s2mPipe_payload_txnId;
      ltAry_5_io_lkResp_s2mPipe_rData_lkType <= ltAry_5_io_lkResp_s2mPipe_payload_lkType;
      ltAry_5_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_5_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_5_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_5_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_5_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_5_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_5_io_lkResp_s2mPipe_rData_wLen <= ltAry_5_io_lkResp_s2mPipe_payload_wLen;
      ltAry_5_io_lkResp_s2mPipe_rData_respType <= ltAry_5_io_lkResp_s2mPipe_payload_respType;
      ltAry_5_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_5_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_6_io_lkResp_ready) begin
      ltAry_6_io_lkResp_rData_nId <= ltAry_6_io_lkResp_payload_nId;
      ltAry_6_io_lkResp_rData_tId <= ltAry_6_io_lkResp_payload_tId;
      ltAry_6_io_lkResp_rData_tabId <= ltAry_6_io_lkResp_payload_tabId;
      ltAry_6_io_lkResp_rData_snId <= ltAry_6_io_lkResp_payload_snId;
      ltAry_6_io_lkResp_rData_txnId <= ltAry_6_io_lkResp_payload_txnId;
      ltAry_6_io_lkResp_rData_lkType <= ltAry_6_io_lkResp_payload_lkType;
      ltAry_6_io_lkResp_rData_lkRelease <= ltAry_6_io_lkResp_payload_lkRelease;
      ltAry_6_io_lkResp_rData_txnAbt <= ltAry_6_io_lkResp_payload_txnAbt;
      ltAry_6_io_lkResp_rData_lkIdx <= ltAry_6_io_lkResp_payload_lkIdx;
      ltAry_6_io_lkResp_rData_wLen <= ltAry_6_io_lkResp_payload_wLen;
      ltAry_6_io_lkResp_rData_respType <= ltAry_6_io_lkResp_payload_respType;
      ltAry_6_io_lkResp_rData_lkWaited <= ltAry_6_io_lkResp_payload_lkWaited;
    end
    if(ltAry_6_io_lkResp_s2mPipe_ready) begin
      ltAry_6_io_lkResp_s2mPipe_rData_nId <= ltAry_6_io_lkResp_s2mPipe_payload_nId;
      ltAry_6_io_lkResp_s2mPipe_rData_tId <= ltAry_6_io_lkResp_s2mPipe_payload_tId;
      ltAry_6_io_lkResp_s2mPipe_rData_tabId <= ltAry_6_io_lkResp_s2mPipe_payload_tabId;
      ltAry_6_io_lkResp_s2mPipe_rData_snId <= ltAry_6_io_lkResp_s2mPipe_payload_snId;
      ltAry_6_io_lkResp_s2mPipe_rData_txnId <= ltAry_6_io_lkResp_s2mPipe_payload_txnId;
      ltAry_6_io_lkResp_s2mPipe_rData_lkType <= ltAry_6_io_lkResp_s2mPipe_payload_lkType;
      ltAry_6_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_6_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_6_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_6_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_6_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_6_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_6_io_lkResp_s2mPipe_rData_wLen <= ltAry_6_io_lkResp_s2mPipe_payload_wLen;
      ltAry_6_io_lkResp_s2mPipe_rData_respType <= ltAry_6_io_lkResp_s2mPipe_payload_respType;
      ltAry_6_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_6_io_lkResp_s2mPipe_payload_lkWaited;
    end
    if(ltAry_7_io_lkResp_ready) begin
      ltAry_7_io_lkResp_rData_nId <= ltAry_7_io_lkResp_payload_nId;
      ltAry_7_io_lkResp_rData_tId <= ltAry_7_io_lkResp_payload_tId;
      ltAry_7_io_lkResp_rData_tabId <= ltAry_7_io_lkResp_payload_tabId;
      ltAry_7_io_lkResp_rData_snId <= ltAry_7_io_lkResp_payload_snId;
      ltAry_7_io_lkResp_rData_txnId <= ltAry_7_io_lkResp_payload_txnId;
      ltAry_7_io_lkResp_rData_lkType <= ltAry_7_io_lkResp_payload_lkType;
      ltAry_7_io_lkResp_rData_lkRelease <= ltAry_7_io_lkResp_payload_lkRelease;
      ltAry_7_io_lkResp_rData_txnAbt <= ltAry_7_io_lkResp_payload_txnAbt;
      ltAry_7_io_lkResp_rData_lkIdx <= ltAry_7_io_lkResp_payload_lkIdx;
      ltAry_7_io_lkResp_rData_wLen <= ltAry_7_io_lkResp_payload_wLen;
      ltAry_7_io_lkResp_rData_respType <= ltAry_7_io_lkResp_payload_respType;
      ltAry_7_io_lkResp_rData_lkWaited <= ltAry_7_io_lkResp_payload_lkWaited;
    end
    if(ltAry_7_io_lkResp_s2mPipe_ready) begin
      ltAry_7_io_lkResp_s2mPipe_rData_nId <= ltAry_7_io_lkResp_s2mPipe_payload_nId;
      ltAry_7_io_lkResp_s2mPipe_rData_tId <= ltAry_7_io_lkResp_s2mPipe_payload_tId;
      ltAry_7_io_lkResp_s2mPipe_rData_tabId <= ltAry_7_io_lkResp_s2mPipe_payload_tabId;
      ltAry_7_io_lkResp_s2mPipe_rData_snId <= ltAry_7_io_lkResp_s2mPipe_payload_snId;
      ltAry_7_io_lkResp_s2mPipe_rData_txnId <= ltAry_7_io_lkResp_s2mPipe_payload_txnId;
      ltAry_7_io_lkResp_s2mPipe_rData_lkType <= ltAry_7_io_lkResp_s2mPipe_payload_lkType;
      ltAry_7_io_lkResp_s2mPipe_rData_lkRelease <= ltAry_7_io_lkResp_s2mPipe_payload_lkRelease;
      ltAry_7_io_lkResp_s2mPipe_rData_txnAbt <= ltAry_7_io_lkResp_s2mPipe_payload_txnAbt;
      ltAry_7_io_lkResp_s2mPipe_rData_lkIdx <= ltAry_7_io_lkResp_s2mPipe_payload_lkIdx;
      ltAry_7_io_lkResp_s2mPipe_rData_wLen <= ltAry_7_io_lkResp_s2mPipe_payload_wLen;
      ltAry_7_io_lkResp_s2mPipe_rData_respType <= ltAry_7_io_lkResp_s2mPipe_payload_respType;
      ltAry_7_io_lkResp_s2mPipe_rData_lkWaited <= ltAry_7_io_lkResp_s2mPipe_payload_lkWaited;
    end
  end


endmodule

//StreamArbiter_5 replaced by StreamArbiter_5

module StreamArbiter_5 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [0:0]    io_inputs_0_payload_nId,
  input      [21:0]   io_inputs_0_payload_tId,
  input      [2:0]    io_inputs_0_payload_tabId,
  input      [0:0]    io_inputs_0_payload_snId,
  input      [5:0]    io_inputs_0_payload_txnId,
  input      [1:0]    io_inputs_0_payload_lkType,
  input               io_inputs_0_payload_lkRelease,
  input               io_inputs_0_payload_txnTimeOut,
  input               io_inputs_0_payload_txnAbt,
  input      [5:0]    io_inputs_0_payload_lkIdx,
  input      [2:0]    io_inputs_0_payload_wLen,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [0:0]    io_inputs_1_payload_nId,
  input      [21:0]   io_inputs_1_payload_tId,
  input      [2:0]    io_inputs_1_payload_tabId,
  input      [0:0]    io_inputs_1_payload_snId,
  input      [5:0]    io_inputs_1_payload_txnId,
  input      [1:0]    io_inputs_1_payload_lkType,
  input               io_inputs_1_payload_lkRelease,
  input               io_inputs_1_payload_txnTimeOut,
  input               io_inputs_1_payload_txnAbt,
  input      [5:0]    io_inputs_1_payload_lkIdx,
  input      [2:0]    io_inputs_1_payload_wLen,
  output              io_output_valid,
  input               io_output_ready,
  output     [0:0]    io_output_payload_nId,
  output     [21:0]   io_output_payload_tId,
  output     [2:0]    io_output_payload_tabId,
  output     [0:0]    io_output_payload_snId,
  output     [5:0]    io_output_payload_txnId,
  output     [1:0]    io_output_payload_lkType,
  output              io_output_payload_lkRelease,
  output              io_output_payload_txnTimeOut,
  output              io_output_payload_txnAbt,
  output     [5:0]    io_output_payload_lkIdx,
  output     [2:0]    io_output_payload_wLen,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire       [1:0]    _zz_io_output_payload_lkType;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [47:0] io_inputs_0_payload_lkType_string;
  reg [47:0] io_inputs_1_payload_lkType_string;
  reg [47:0] io_output_payload_lkType_string;
  reg [47:0] _zz_io_output_payload_lkType_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_lkType)
      LkT_rd : io_inputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_0_payload_lkType_string = "insTab";
      default : io_inputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_lkType)
      LkT_rd : io_inputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_1_payload_lkType_string = "insTab";
      default : io_inputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_lkType)
      LkT_rd : io_output_payload_lkType_string = "rd    ";
      LkT_wr : io_output_payload_lkType_string = "wr    ";
      LkT_raw : io_output_payload_lkType_string = "raw   ";
      LkT_insTab : io_output_payload_lkType_string = "insTab";
      default : io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_lkType)
      LkT_rd : _zz_io_output_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_output_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_output_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_output_payload_lkType_string = "insTab";
      default : _zz_io_output_payload_lkType_string = "??????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_lkType = (maskRouted_0 ? io_inputs_0_payload_lkType : io_inputs_1_payload_lkType);
  assign io_output_payload_nId = (maskRouted_0 ? io_inputs_0_payload_nId : io_inputs_1_payload_nId);
  assign io_output_payload_tId = (maskRouted_0 ? io_inputs_0_payload_tId : io_inputs_1_payload_tId);
  assign io_output_payload_tabId = (maskRouted_0 ? io_inputs_0_payload_tabId : io_inputs_1_payload_tabId);
  assign io_output_payload_snId = (maskRouted_0 ? io_inputs_0_payload_snId : io_inputs_1_payload_snId);
  assign io_output_payload_txnId = (maskRouted_0 ? io_inputs_0_payload_txnId : io_inputs_1_payload_txnId);
  assign io_output_payload_lkType = _zz_io_output_payload_lkType;
  assign io_output_payload_lkRelease = (maskRouted_0 ? io_inputs_0_payload_lkRelease : io_inputs_1_payload_lkRelease);
  assign io_output_payload_txnTimeOut = (maskRouted_0 ? io_inputs_0_payload_txnTimeOut : io_inputs_1_payload_txnTimeOut);
  assign io_output_payload_txnAbt = (maskRouted_0 ? io_inputs_0_payload_txnAbt : io_inputs_1_payload_txnAbt);
  assign io_output_payload_lkIdx = (maskRouted_0 ? io_inputs_0_payload_lkIdx : io_inputs_1_payload_lkIdx);
  assign io_output_payload_wLen = (maskRouted_0 ? io_inputs_0_payload_wLen : io_inputs_1_payload_wLen);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(!resetn) begin
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
    end
  end


endmodule

//StreamArbiter_3 replaced by StreamArbiter_3

module StreamArbiter_3 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [0:0]    io_inputs_0_payload_nId,
  input      [21:0]   io_inputs_0_payload_tId,
  input      [2:0]    io_inputs_0_payload_tabId,
  input      [0:0]    io_inputs_0_payload_snId,
  input      [5:0]    io_inputs_0_payload_txnId,
  input      [1:0]    io_inputs_0_payload_lkType,
  input               io_inputs_0_payload_lkRelease,
  input               io_inputs_0_payload_txnAbt,
  input      [5:0]    io_inputs_0_payload_lkIdx,
  input      [2:0]    io_inputs_0_payload_wLen,
  input      [1:0]    io_inputs_0_payload_respType,
  input               io_inputs_0_payload_lkWaited,
  output              io_output_valid,
  input               io_output_ready,
  output     [0:0]    io_output_payload_nId,
  output     [21:0]   io_output_payload_tId,
  output     [2:0]    io_output_payload_tabId,
  output     [0:0]    io_output_payload_snId,
  output     [5:0]    io_output_payload_txnId,
  output     [1:0]    io_output_payload_lkType,
  output              io_output_payload_lkRelease,
  output              io_output_payload_txnAbt,
  output     [5:0]    io_output_payload_lkIdx,
  output     [2:0]    io_output_payload_wLen,
  output     [1:0]    io_output_payload_respType,
  output              io_output_payload_lkWaited,
  output     [0:0]    io_chosenOH,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire       [1:0]    _zz__zz_maskProposal_0_2;
  wire       [1:0]    _zz__zz_maskProposal_0_2_1;
  wire       [0:0]    _zz__zz_maskProposal_0_2_2;
  wire       [0:0]    _zz_maskProposal_0_3;
  reg                 locked;
  wire                maskProposal_0;
  reg                 maskLocked_0;
  wire                maskRouted_0;
  wire       [0:0]    _zz_maskProposal_0;
  wire       [1:0]    _zz_maskProposal_0_1;
  wire       [1:0]    _zz_maskProposal_0_2;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_lkType;
  wire       [1:0]    _zz_io_output_payload_respType;
  `ifndef SYNTHESIS
  reg [47:0] io_inputs_0_payload_lkType_string;
  reg [71:0] io_inputs_0_payload_respType_string;
  reg [47:0] io_output_payload_lkType_string;
  reg [71:0] io_output_payload_respType_string;
  reg [47:0] _zz_io_output_payload_lkType_string;
  reg [71:0] _zz_io_output_payload_respType_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = maskLocked_0;
  assign _zz__zz_maskProposal_0_2_1 = {1'd0, _zz__zz_maskProposal_0_2_2};
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[1 : 1] | _zz_maskProposal_0_2[0 : 0]);
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_lkType)
      LkT_rd : io_inputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_0_payload_lkType_string = "insTab";
      default : io_inputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_respType)
      LockRespType_grant : io_inputs_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_0_payload_respType_string = "release_1";
      default : io_inputs_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_lkType)
      LkT_rd : io_output_payload_lkType_string = "rd    ";
      LkT_wr : io_output_payload_lkType_string = "wr    ";
      LkT_raw : io_output_payload_lkType_string = "raw   ";
      LkT_insTab : io_output_payload_lkType_string = "insTab";
      default : io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_respType)
      LockRespType_grant : io_output_payload_respType_string = "grant    ";
      LockRespType_abort : io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_output_payload_respType_string = "release_1";
      default : io_output_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_lkType)
      LkT_rd : _zz_io_output_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_output_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_output_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_output_payload_lkType_string = "insTab";
      default : _zz_io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_respType)
      LockRespType_grant : _zz_io_output_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_io_output_payload_respType_string = "release_1";
      default : _zz_io_output_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign _zz_maskProposal_0 = io_inputs_0_valid;
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (io_inputs_0_valid && maskRouted_0);
  assign _zz_io_output_payload_lkType = io_inputs_0_payload_lkType;
  assign _zz_io_output_payload_respType = io_inputs_0_payload_respType;
  assign io_output_payload_nId = io_inputs_0_payload_nId;
  assign io_output_payload_tId = io_inputs_0_payload_tId;
  assign io_output_payload_tabId = io_inputs_0_payload_tabId;
  assign io_output_payload_snId = io_inputs_0_payload_snId;
  assign io_output_payload_txnId = io_inputs_0_payload_txnId;
  assign io_output_payload_lkType = _zz_io_output_payload_lkType;
  assign io_output_payload_lkRelease = io_inputs_0_payload_lkRelease;
  assign io_output_payload_txnAbt = io_inputs_0_payload_txnAbt;
  assign io_output_payload_lkIdx = io_inputs_0_payload_lkIdx;
  assign io_output_payload_wLen = io_inputs_0_payload_wLen;
  assign io_output_payload_respType = _zz_io_output_payload_respType;
  assign io_output_payload_lkWaited = io_inputs_0_payload_lkWaited;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_chosenOH = maskRouted_0;
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamDemux2_2 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [0:0]    io_input_payload_nId,
  input      [21:0]   io_input_payload_tId,
  input      [2:0]    io_input_payload_tabId,
  input      [0:0]    io_input_payload_snId,
  input      [5:0]    io_input_payload_txnId,
  input      [1:0]    io_input_payload_lkType,
  input               io_input_payload_lkRelease,
  input               io_input_payload_txnAbt,
  input      [5:0]    io_input_payload_lkIdx,
  input      [2:0]    io_input_payload_wLen,
  input      [1:0]    io_input_payload_respType,
  input               io_input_payload_lkWaited,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [0:0]    io_outputs_0_payload_nId,
  output     [21:0]   io_outputs_0_payload_tId,
  output     [2:0]    io_outputs_0_payload_tabId,
  output     [0:0]    io_outputs_0_payload_snId,
  output     [5:0]    io_outputs_0_payload_txnId,
  output     [1:0]    io_outputs_0_payload_lkType,
  output              io_outputs_0_payload_lkRelease,
  output              io_outputs_0_payload_txnAbt,
  output     [5:0]    io_outputs_0_payload_lkIdx,
  output     [2:0]    io_outputs_0_payload_wLen,
  output     [1:0]    io_outputs_0_payload_respType,
  output              io_outputs_0_payload_lkWaited,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [0:0]    io_outputs_1_payload_nId,
  output     [21:0]   io_outputs_1_payload_tId,
  output     [2:0]    io_outputs_1_payload_tabId,
  output     [0:0]    io_outputs_1_payload_snId,
  output     [5:0]    io_outputs_1_payload_txnId,
  output     [1:0]    io_outputs_1_payload_lkType,
  output              io_outputs_1_payload_lkRelease,
  output              io_outputs_1_payload_txnAbt,
  output     [5:0]    io_outputs_1_payload_lkIdx,
  output     [2:0]    io_outputs_1_payload_wLen,
  output     [1:0]    io_outputs_1_payload_respType,
  output              io_outputs_1_payload_lkWaited
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire                when_Interconnect_l54;
  wire                when_Interconnect_l54_1;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_lkType_string;
  reg [71:0] io_input_payload_respType_string;
  reg [47:0] io_outputs_0_payload_lkType_string;
  reg [71:0] io_outputs_0_payload_respType_string;
  reg [47:0] io_outputs_1_payload_lkType_string;
  reg [71:0] io_outputs_1_payload_respType_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_lkType)
      LkT_rd : io_input_payload_lkType_string = "rd    ";
      LkT_wr : io_input_payload_lkType_string = "wr    ";
      LkT_raw : io_input_payload_lkType_string = "raw   ";
      LkT_insTab : io_input_payload_lkType_string = "insTab";
      default : io_input_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_input_payload_respType)
      LockRespType_grant : io_input_payload_respType_string = "grant    ";
      LockRespType_abort : io_input_payload_respType_string = "abort    ";
      LockRespType_waiting : io_input_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_input_payload_respType_string = "release_1";
      default : io_input_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_lkType)
      LkT_rd : io_outputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_0_payload_lkType_string = "insTab";
      default : io_outputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_respType)
      LockRespType_grant : io_outputs_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_outputs_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_outputs_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_outputs_0_payload_respType_string = "release_1";
      default : io_outputs_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_lkType)
      LkT_rd : io_outputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_1_payload_lkType_string = "insTab";
      default : io_outputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_respType)
      LockRespType_grant : io_outputs_1_payload_respType_string = "grant    ";
      LockRespType_abort : io_outputs_1_payload_respType_string = "abort    ";
      LockRespType_waiting : io_outputs_1_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_outputs_1_payload_respType_string = "release_1";
      default : io_outputs_1_payload_respType_string = "?????????";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Interconnect_l54) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Interconnect_l54_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_nId = io_input_payload_nId;
  assign io_outputs_0_payload_tId = io_input_payload_tId;
  assign io_outputs_0_payload_tabId = io_input_payload_tabId;
  assign io_outputs_0_payload_snId = io_input_payload_snId;
  assign io_outputs_0_payload_txnId = io_input_payload_txnId;
  assign io_outputs_0_payload_lkType = io_input_payload_lkType;
  assign io_outputs_0_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_0_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_0_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_0_payload_wLen = io_input_payload_wLen;
  assign io_outputs_0_payload_respType = io_input_payload_respType;
  assign io_outputs_0_payload_lkWaited = io_input_payload_lkWaited;
  assign when_Interconnect_l54 = (1'b0 != io_select);
  always @(*) begin
    if(when_Interconnect_l54) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_nId = io_input_payload_nId;
  assign io_outputs_1_payload_tId = io_input_payload_tId;
  assign io_outputs_1_payload_tabId = io_input_payload_tabId;
  assign io_outputs_1_payload_snId = io_input_payload_snId;
  assign io_outputs_1_payload_txnId = io_input_payload_txnId;
  assign io_outputs_1_payload_lkType = io_input_payload_lkType;
  assign io_outputs_1_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_1_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_1_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_1_payload_wLen = io_input_payload_wLen;
  assign io_outputs_1_payload_respType = io_input_payload_respType;
  assign io_outputs_1_payload_lkWaited = io_input_payload_lkWaited;
  assign when_Interconnect_l54_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Interconnect_l54_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module StreamArbiter_2 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [0:0]    io_inputs_0_payload_nId,
  input      [21:0]   io_inputs_0_payload_tId,
  input      [2:0]    io_inputs_0_payload_tabId,
  input      [0:0]    io_inputs_0_payload_snId,
  input      [5:0]    io_inputs_0_payload_txnId,
  input      [1:0]    io_inputs_0_payload_lkType,
  input               io_inputs_0_payload_lkRelease,
  input               io_inputs_0_payload_txnTimeOut,
  input               io_inputs_0_payload_txnAbt,
  input      [5:0]    io_inputs_0_payload_lkIdx,
  input      [2:0]    io_inputs_0_payload_wLen,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [0:0]    io_inputs_1_payload_nId,
  input      [21:0]   io_inputs_1_payload_tId,
  input      [2:0]    io_inputs_1_payload_tabId,
  input      [0:0]    io_inputs_1_payload_snId,
  input      [5:0]    io_inputs_1_payload_txnId,
  input      [1:0]    io_inputs_1_payload_lkType,
  input               io_inputs_1_payload_lkRelease,
  input               io_inputs_1_payload_txnTimeOut,
  input               io_inputs_1_payload_txnAbt,
  input      [5:0]    io_inputs_1_payload_lkIdx,
  input      [2:0]    io_inputs_1_payload_wLen,
  output              io_output_valid,
  input               io_output_ready,
  output     [0:0]    io_output_payload_nId,
  output     [21:0]   io_output_payload_tId,
  output     [2:0]    io_output_payload_tabId,
  output     [0:0]    io_output_payload_snId,
  output     [5:0]    io_output_payload_txnId,
  output     [1:0]    io_output_payload_lkType,
  output              io_output_payload_lkRelease,
  output              io_output_payload_txnTimeOut,
  output              io_output_payload_txnAbt,
  output     [5:0]    io_output_payload_lkIdx,
  output     [2:0]    io_output_payload_wLen,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_lkType;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [47:0] io_inputs_0_payload_lkType_string;
  reg [47:0] io_inputs_1_payload_lkType_string;
  reg [47:0] io_output_payload_lkType_string;
  reg [47:0] _zz_io_output_payload_lkType_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_lkType)
      LkT_rd : io_inputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_0_payload_lkType_string = "insTab";
      default : io_inputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_lkType)
      LkT_rd : io_inputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_1_payload_lkType_string = "insTab";
      default : io_inputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_lkType)
      LkT_rd : io_output_payload_lkType_string = "rd    ";
      LkT_wr : io_output_payload_lkType_string = "wr    ";
      LkT_raw : io_output_payload_lkType_string = "raw   ";
      LkT_insTab : io_output_payload_lkType_string = "insTab";
      default : io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_lkType)
      LkT_rd : _zz_io_output_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_output_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_output_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_output_payload_lkType_string = "insTab";
      default : _zz_io_output_payload_lkType_string = "??????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_lkType = (maskRouted_0 ? io_inputs_0_payload_lkType : io_inputs_1_payload_lkType);
  assign io_output_payload_nId = (maskRouted_0 ? io_inputs_0_payload_nId : io_inputs_1_payload_nId);
  assign io_output_payload_tId = (maskRouted_0 ? io_inputs_0_payload_tId : io_inputs_1_payload_tId);
  assign io_output_payload_tabId = (maskRouted_0 ? io_inputs_0_payload_tabId : io_inputs_1_payload_tabId);
  assign io_output_payload_snId = (maskRouted_0 ? io_inputs_0_payload_snId : io_inputs_1_payload_snId);
  assign io_output_payload_txnId = (maskRouted_0 ? io_inputs_0_payload_txnId : io_inputs_1_payload_txnId);
  assign io_output_payload_lkType = _zz_io_output_payload_lkType;
  assign io_output_payload_lkRelease = (maskRouted_0 ? io_inputs_0_payload_lkRelease : io_inputs_1_payload_lkRelease);
  assign io_output_payload_txnTimeOut = (maskRouted_0 ? io_inputs_0_payload_txnTimeOut : io_inputs_1_payload_txnTimeOut);
  assign io_output_payload_txnAbt = (maskRouted_0 ? io_inputs_0_payload_txnAbt : io_inputs_1_payload_txnAbt);
  assign io_output_payload_lkIdx = (maskRouted_0 ? io_inputs_0_payload_lkIdx : io_inputs_1_payload_lkIdx);
  assign io_output_payload_wLen = (maskRouted_0 ? io_inputs_0_payload_wLen : io_inputs_1_payload_wLen);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

//StreamDemux2 replaced by StreamDemux2

module StreamDemux2 (
  input               io_input_valid,
  output reg          io_input_ready,
  input      [0:0]    io_input_payload_nId,
  input      [21:0]   io_input_payload_tId,
  input      [2:0]    io_input_payload_tabId,
  input      [0:0]    io_input_payload_snId,
  input      [5:0]    io_input_payload_txnId,
  input      [1:0]    io_input_payload_lkType,
  input               io_input_payload_lkRelease,
  input               io_input_payload_txnTimeOut,
  input               io_input_payload_txnAbt,
  input      [5:0]    io_input_payload_lkIdx,
  input      [2:0]    io_input_payload_wLen,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [0:0]    io_outputs_0_payload_nId,
  output     [21:0]   io_outputs_0_payload_tId,
  output     [2:0]    io_outputs_0_payload_tabId,
  output     [0:0]    io_outputs_0_payload_snId,
  output     [5:0]    io_outputs_0_payload_txnId,
  output     [1:0]    io_outputs_0_payload_lkType,
  output              io_outputs_0_payload_lkRelease,
  output              io_outputs_0_payload_txnTimeOut,
  output              io_outputs_0_payload_txnAbt,
  output     [5:0]    io_outputs_0_payload_lkIdx,
  output     [2:0]    io_outputs_0_payload_wLen
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire                when_Interconnect_l54;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_lkType_string;
  reg [47:0] io_outputs_0_payload_lkType_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_lkType)
      LkT_rd : io_input_payload_lkType_string = "rd    ";
      LkT_wr : io_input_payload_lkType_string = "wr    ";
      LkT_raw : io_input_payload_lkType_string = "raw   ";
      LkT_insTab : io_input_payload_lkType_string = "insTab";
      default : io_input_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_lkType)
      LkT_rd : io_outputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_0_payload_lkType_string = "insTab";
      default : io_outputs_0_payload_lkType_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Interconnect_l54) begin
      io_input_ready = io_outputs_0_ready;
    end
  end

  assign io_outputs_0_payload_nId = io_input_payload_nId;
  assign io_outputs_0_payload_tId = io_input_payload_tId;
  assign io_outputs_0_payload_tabId = io_input_payload_tabId;
  assign io_outputs_0_payload_snId = io_input_payload_snId;
  assign io_outputs_0_payload_txnId = io_input_payload_txnId;
  assign io_outputs_0_payload_lkType = io_input_payload_lkType;
  assign io_outputs_0_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_0_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_0_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_0_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_0_payload_wLen = io_input_payload_wLen;
  assign when_Interconnect_l54 = 1'b0;
  always @(*) begin
    if(when_Interconnect_l54) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end


endmodule

module StreamArbiter_1 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [0:0]    io_inputs_0_payload_nId,
  input      [21:0]   io_inputs_0_payload_tId,
  input      [2:0]    io_inputs_0_payload_tabId,
  input      [0:0]    io_inputs_0_payload_snId,
  input      [5:0]    io_inputs_0_payload_txnId,
  input      [1:0]    io_inputs_0_payload_lkType,
  input               io_inputs_0_payload_lkRelease,
  input               io_inputs_0_payload_txnAbt,
  input      [5:0]    io_inputs_0_payload_lkIdx,
  input      [2:0]    io_inputs_0_payload_wLen,
  input      [1:0]    io_inputs_0_payload_respType,
  input               io_inputs_0_payload_lkWaited,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [0:0]    io_inputs_1_payload_nId,
  input      [21:0]   io_inputs_1_payload_tId,
  input      [2:0]    io_inputs_1_payload_tabId,
  input      [0:0]    io_inputs_1_payload_snId,
  input      [5:0]    io_inputs_1_payload_txnId,
  input      [1:0]    io_inputs_1_payload_lkType,
  input               io_inputs_1_payload_lkRelease,
  input               io_inputs_1_payload_txnAbt,
  input      [5:0]    io_inputs_1_payload_lkIdx,
  input      [2:0]    io_inputs_1_payload_wLen,
  input      [1:0]    io_inputs_1_payload_respType,
  input               io_inputs_1_payload_lkWaited,
  output              io_output_valid,
  input               io_output_ready,
  output     [0:0]    io_output_payload_nId,
  output     [21:0]   io_output_payload_tId,
  output     [2:0]    io_output_payload_tabId,
  output     [0:0]    io_output_payload_snId,
  output     [5:0]    io_output_payload_txnId,
  output     [1:0]    io_output_payload_lkType,
  output              io_output_payload_lkRelease,
  output              io_output_payload_txnAbt,
  output     [5:0]    io_output_payload_lkIdx,
  output     [2:0]    io_output_payload_wLen,
  output     [1:0]    io_output_payload_respType,
  output              io_output_payload_lkWaited,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_lkType;
  wire       [1:0]    _zz_io_output_payload_respType;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [47:0] io_inputs_0_payload_lkType_string;
  reg [71:0] io_inputs_0_payload_respType_string;
  reg [47:0] io_inputs_1_payload_lkType_string;
  reg [71:0] io_inputs_1_payload_respType_string;
  reg [47:0] io_output_payload_lkType_string;
  reg [71:0] io_output_payload_respType_string;
  reg [47:0] _zz_io_output_payload_lkType_string;
  reg [71:0] _zz_io_output_payload_respType_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_lkType)
      LkT_rd : io_inputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_0_payload_lkType_string = "insTab";
      default : io_inputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_respType)
      LockRespType_grant : io_inputs_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_0_payload_respType_string = "release_1";
      default : io_inputs_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_lkType)
      LkT_rd : io_inputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_1_payload_lkType_string = "insTab";
      default : io_inputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_respType)
      LockRespType_grant : io_inputs_1_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_1_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_1_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_1_payload_respType_string = "release_1";
      default : io_inputs_1_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_lkType)
      LkT_rd : io_output_payload_lkType_string = "rd    ";
      LkT_wr : io_output_payload_lkType_string = "wr    ";
      LkT_raw : io_output_payload_lkType_string = "raw   ";
      LkT_insTab : io_output_payload_lkType_string = "insTab";
      default : io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_respType)
      LockRespType_grant : io_output_payload_respType_string = "grant    ";
      LockRespType_abort : io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_output_payload_respType_string = "release_1";
      default : io_output_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_lkType)
      LkT_rd : _zz_io_output_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_output_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_output_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_output_payload_lkType_string = "insTab";
      default : _zz_io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_respType)
      LockRespType_grant : _zz_io_output_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_io_output_payload_respType_string = "release_1";
      default : _zz_io_output_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_lkType = (maskRouted_0 ? io_inputs_0_payload_lkType : io_inputs_1_payload_lkType);
  assign _zz_io_output_payload_respType = (maskRouted_0 ? io_inputs_0_payload_respType : io_inputs_1_payload_respType);
  assign io_output_payload_nId = (maskRouted_0 ? io_inputs_0_payload_nId : io_inputs_1_payload_nId);
  assign io_output_payload_tId = (maskRouted_0 ? io_inputs_0_payload_tId : io_inputs_1_payload_tId);
  assign io_output_payload_tabId = (maskRouted_0 ? io_inputs_0_payload_tabId : io_inputs_1_payload_tabId);
  assign io_output_payload_snId = (maskRouted_0 ? io_inputs_0_payload_snId : io_inputs_1_payload_snId);
  assign io_output_payload_txnId = (maskRouted_0 ? io_inputs_0_payload_txnId : io_inputs_1_payload_txnId);
  assign io_output_payload_lkType = _zz_io_output_payload_lkType;
  assign io_output_payload_lkRelease = (maskRouted_0 ? io_inputs_0_payload_lkRelease : io_inputs_1_payload_lkRelease);
  assign io_output_payload_txnAbt = (maskRouted_0 ? io_inputs_0_payload_txnAbt : io_inputs_1_payload_txnAbt);
  assign io_output_payload_lkIdx = (maskRouted_0 ? io_inputs_0_payload_lkIdx : io_inputs_1_payload_lkIdx);
  assign io_output_payload_wLen = (maskRouted_0 ? io_inputs_0_payload_wLen : io_inputs_1_payload_wLen);
  assign io_output_payload_respType = _zz_io_output_payload_respType;
  assign io_output_payload_lkWaited = (maskRouted_0 ? io_inputs_0_payload_lkWaited : io_inputs_1_payload_lkWaited);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [0:0]    io_inputs_0_payload_nId,
  input      [18:0]   io_inputs_0_payload_tId,
  input      [2:0]    io_inputs_0_payload_tabId,
  input      [0:0]    io_inputs_0_payload_snId,
  input      [5:0]    io_inputs_0_payload_txnId,
  input      [1:0]    io_inputs_0_payload_lkType,
  input               io_inputs_0_payload_lkRelease,
  input               io_inputs_0_payload_txnAbt,
  input      [5:0]    io_inputs_0_payload_lkIdx,
  input      [2:0]    io_inputs_0_payload_wLen,
  input      [1:0]    io_inputs_0_payload_respType,
  input               io_inputs_0_payload_lkWaited,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [0:0]    io_inputs_1_payload_nId,
  input      [18:0]   io_inputs_1_payload_tId,
  input      [2:0]    io_inputs_1_payload_tabId,
  input      [0:0]    io_inputs_1_payload_snId,
  input      [5:0]    io_inputs_1_payload_txnId,
  input      [1:0]    io_inputs_1_payload_lkType,
  input               io_inputs_1_payload_lkRelease,
  input               io_inputs_1_payload_txnAbt,
  input      [5:0]    io_inputs_1_payload_lkIdx,
  input      [2:0]    io_inputs_1_payload_wLen,
  input      [1:0]    io_inputs_1_payload_respType,
  input               io_inputs_1_payload_lkWaited,
  input               io_inputs_2_valid,
  output              io_inputs_2_ready,
  input      [0:0]    io_inputs_2_payload_nId,
  input      [18:0]   io_inputs_2_payload_tId,
  input      [2:0]    io_inputs_2_payload_tabId,
  input      [0:0]    io_inputs_2_payload_snId,
  input      [5:0]    io_inputs_2_payload_txnId,
  input      [1:0]    io_inputs_2_payload_lkType,
  input               io_inputs_2_payload_lkRelease,
  input               io_inputs_2_payload_txnAbt,
  input      [5:0]    io_inputs_2_payload_lkIdx,
  input      [2:0]    io_inputs_2_payload_wLen,
  input      [1:0]    io_inputs_2_payload_respType,
  input               io_inputs_2_payload_lkWaited,
  input               io_inputs_3_valid,
  output              io_inputs_3_ready,
  input      [0:0]    io_inputs_3_payload_nId,
  input      [18:0]   io_inputs_3_payload_tId,
  input      [2:0]    io_inputs_3_payload_tabId,
  input      [0:0]    io_inputs_3_payload_snId,
  input      [5:0]    io_inputs_3_payload_txnId,
  input      [1:0]    io_inputs_3_payload_lkType,
  input               io_inputs_3_payload_lkRelease,
  input               io_inputs_3_payload_txnAbt,
  input      [5:0]    io_inputs_3_payload_lkIdx,
  input      [2:0]    io_inputs_3_payload_wLen,
  input      [1:0]    io_inputs_3_payload_respType,
  input               io_inputs_3_payload_lkWaited,
  input               io_inputs_4_valid,
  output              io_inputs_4_ready,
  input      [0:0]    io_inputs_4_payload_nId,
  input      [18:0]   io_inputs_4_payload_tId,
  input      [2:0]    io_inputs_4_payload_tabId,
  input      [0:0]    io_inputs_4_payload_snId,
  input      [5:0]    io_inputs_4_payload_txnId,
  input      [1:0]    io_inputs_4_payload_lkType,
  input               io_inputs_4_payload_lkRelease,
  input               io_inputs_4_payload_txnAbt,
  input      [5:0]    io_inputs_4_payload_lkIdx,
  input      [2:0]    io_inputs_4_payload_wLen,
  input      [1:0]    io_inputs_4_payload_respType,
  input               io_inputs_4_payload_lkWaited,
  input               io_inputs_5_valid,
  output              io_inputs_5_ready,
  input      [0:0]    io_inputs_5_payload_nId,
  input      [18:0]   io_inputs_5_payload_tId,
  input      [2:0]    io_inputs_5_payload_tabId,
  input      [0:0]    io_inputs_5_payload_snId,
  input      [5:0]    io_inputs_5_payload_txnId,
  input      [1:0]    io_inputs_5_payload_lkType,
  input               io_inputs_5_payload_lkRelease,
  input               io_inputs_5_payload_txnAbt,
  input      [5:0]    io_inputs_5_payload_lkIdx,
  input      [2:0]    io_inputs_5_payload_wLen,
  input      [1:0]    io_inputs_5_payload_respType,
  input               io_inputs_5_payload_lkWaited,
  input               io_inputs_6_valid,
  output              io_inputs_6_ready,
  input      [0:0]    io_inputs_6_payload_nId,
  input      [18:0]   io_inputs_6_payload_tId,
  input      [2:0]    io_inputs_6_payload_tabId,
  input      [0:0]    io_inputs_6_payload_snId,
  input      [5:0]    io_inputs_6_payload_txnId,
  input      [1:0]    io_inputs_6_payload_lkType,
  input               io_inputs_6_payload_lkRelease,
  input               io_inputs_6_payload_txnAbt,
  input      [5:0]    io_inputs_6_payload_lkIdx,
  input      [2:0]    io_inputs_6_payload_wLen,
  input      [1:0]    io_inputs_6_payload_respType,
  input               io_inputs_6_payload_lkWaited,
  input               io_inputs_7_valid,
  output              io_inputs_7_ready,
  input      [0:0]    io_inputs_7_payload_nId,
  input      [18:0]   io_inputs_7_payload_tId,
  input      [2:0]    io_inputs_7_payload_tabId,
  input      [0:0]    io_inputs_7_payload_snId,
  input      [5:0]    io_inputs_7_payload_txnId,
  input      [1:0]    io_inputs_7_payload_lkType,
  input               io_inputs_7_payload_lkRelease,
  input               io_inputs_7_payload_txnAbt,
  input      [5:0]    io_inputs_7_payload_lkIdx,
  input      [2:0]    io_inputs_7_payload_wLen,
  input      [1:0]    io_inputs_7_payload_respType,
  input               io_inputs_7_payload_lkWaited,
  output              io_output_valid,
  input               io_output_ready,
  output     [0:0]    io_output_payload_nId,
  output     [18:0]   io_output_payload_tId,
  output     [2:0]    io_output_payload_tabId,
  output     [0:0]    io_output_payload_snId,
  output     [5:0]    io_output_payload_txnId,
  output     [1:0]    io_output_payload_lkType,
  output              io_output_payload_lkRelease,
  output              io_output_payload_txnAbt,
  output     [5:0]    io_output_payload_lkIdx,
  output     [2:0]    io_output_payload_wLen,
  output     [1:0]    io_output_payload_respType,
  output              io_output_payload_lkWaited,
  output     [2:0]    io_chosen,
  output     [7:0]    io_chosenOH,
  input               clk,
  input               resetn
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;

  wire       [15:0]   _zz__zz_maskProposal_0_2;
  wire       [15:0]   _zz__zz_maskProposal_0_2_1;
  wire       [7:0]    _zz__zz_maskProposal_0_2_2;
  reg        [1:0]    _zz__zz_io_output_payload_lkType;
  reg        [1:0]    _zz__zz_io_output_payload_respType;
  reg        [0:0]    _zz_io_output_payload_nId_4;
  reg        [18:0]   _zz_io_output_payload_tId;
  reg        [2:0]    _zz_io_output_payload_tabId;
  reg        [0:0]    _zz_io_output_payload_snId;
  reg        [5:0]    _zz_io_output_payload_txnId;
  reg                 _zz_io_output_payload_lkRelease;
  reg                 _zz_io_output_payload_txnAbt;
  reg        [5:0]    _zz_io_output_payload_lkIdx;
  reg        [2:0]    _zz_io_output_payload_wLen;
  reg                 _zz_io_output_payload_lkWaited;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  wire                maskProposal_4;
  wire                maskProposal_5;
  wire                maskProposal_6;
  wire                maskProposal_7;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  reg                 maskLocked_4;
  reg                 maskLocked_5;
  reg                 maskLocked_6;
  reg                 maskLocked_7;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire                maskRouted_4;
  wire                maskRouted_5;
  wire                maskRouted_6;
  wire                maskRouted_7;
  wire       [7:0]    _zz_maskProposal_0;
  wire       [15:0]   _zz_maskProposal_0_1;
  wire       [15:0]   _zz_maskProposal_0_2;
  wire       [7:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_output_payload_nId;
  wire                _zz_io_output_payload_nId_1;
  wire                _zz_io_output_payload_nId_2;
  wire       [2:0]    _zz_io_output_payload_nId_3;
  wire       [1:0]    _zz_io_output_payload_lkType;
  wire       [1:0]    _zz_io_output_payload_respType;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;
  wire                _zz_io_chosen_3;
  wire                _zz_io_chosen_4;
  wire                _zz_io_chosen_5;
  wire                _zz_io_chosen_6;
  `ifndef SYNTHESIS
  reg [47:0] io_inputs_0_payload_lkType_string;
  reg [71:0] io_inputs_0_payload_respType_string;
  reg [47:0] io_inputs_1_payload_lkType_string;
  reg [71:0] io_inputs_1_payload_respType_string;
  reg [47:0] io_inputs_2_payload_lkType_string;
  reg [71:0] io_inputs_2_payload_respType_string;
  reg [47:0] io_inputs_3_payload_lkType_string;
  reg [71:0] io_inputs_3_payload_respType_string;
  reg [47:0] io_inputs_4_payload_lkType_string;
  reg [71:0] io_inputs_4_payload_respType_string;
  reg [47:0] io_inputs_5_payload_lkType_string;
  reg [71:0] io_inputs_5_payload_respType_string;
  reg [47:0] io_inputs_6_payload_lkType_string;
  reg [71:0] io_inputs_6_payload_respType_string;
  reg [47:0] io_inputs_7_payload_lkType_string;
  reg [71:0] io_inputs_7_payload_respType_string;
  reg [47:0] io_output_payload_lkType_string;
  reg [71:0] io_output_payload_respType_string;
  reg [47:0] _zz_io_output_payload_lkType_string;
  reg [71:0] _zz_io_output_payload_respType_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_6,{maskLocked_5,{maskLocked_4,{maskLocked_3,{maskLocked_2,{maskLocked_1,{maskLocked_0,maskLocked_7}}}}}}};
  assign _zz__zz_maskProposal_0_2_1 = {8'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_nId_3)
      3'b000 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_0_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_0_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_0_payload_nId;
        _zz_io_output_payload_tId = io_inputs_0_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_0_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_0_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_0_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_0_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_0_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_0_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_0_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_0_payload_lkWaited;
      end
      3'b001 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_1_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_1_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_1_payload_nId;
        _zz_io_output_payload_tId = io_inputs_1_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_1_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_1_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_1_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_1_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_1_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_1_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_1_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_1_payload_lkWaited;
      end
      3'b010 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_2_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_2_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_2_payload_nId;
        _zz_io_output_payload_tId = io_inputs_2_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_2_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_2_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_2_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_2_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_2_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_2_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_2_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_2_payload_lkWaited;
      end
      3'b011 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_3_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_3_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_3_payload_nId;
        _zz_io_output_payload_tId = io_inputs_3_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_3_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_3_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_3_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_3_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_3_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_3_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_3_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_3_payload_lkWaited;
      end
      3'b100 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_4_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_4_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_4_payload_nId;
        _zz_io_output_payload_tId = io_inputs_4_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_4_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_4_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_4_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_4_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_4_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_4_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_4_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_4_payload_lkWaited;
      end
      3'b101 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_5_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_5_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_5_payload_nId;
        _zz_io_output_payload_tId = io_inputs_5_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_5_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_5_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_5_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_5_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_5_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_5_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_5_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_5_payload_lkWaited;
      end
      3'b110 : begin
        _zz__zz_io_output_payload_lkType = io_inputs_6_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_6_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_6_payload_nId;
        _zz_io_output_payload_tId = io_inputs_6_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_6_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_6_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_6_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_6_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_6_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_6_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_6_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_6_payload_lkWaited;
      end
      default : begin
        _zz__zz_io_output_payload_lkType = io_inputs_7_payload_lkType;
        _zz__zz_io_output_payload_respType = io_inputs_7_payload_respType;
        _zz_io_output_payload_nId_4 = io_inputs_7_payload_nId;
        _zz_io_output_payload_tId = io_inputs_7_payload_tId;
        _zz_io_output_payload_tabId = io_inputs_7_payload_tabId;
        _zz_io_output_payload_snId = io_inputs_7_payload_snId;
        _zz_io_output_payload_txnId = io_inputs_7_payload_txnId;
        _zz_io_output_payload_lkRelease = io_inputs_7_payload_lkRelease;
        _zz_io_output_payload_txnAbt = io_inputs_7_payload_txnAbt;
        _zz_io_output_payload_lkIdx = io_inputs_7_payload_lkIdx;
        _zz_io_output_payload_wLen = io_inputs_7_payload_wLen;
        _zz_io_output_payload_lkWaited = io_inputs_7_payload_lkWaited;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_lkType)
      LkT_rd : io_inputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_0_payload_lkType_string = "insTab";
      default : io_inputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_respType)
      LockRespType_grant : io_inputs_0_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_0_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_0_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_0_payload_respType_string = "release_1";
      default : io_inputs_0_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_lkType)
      LkT_rd : io_inputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_1_payload_lkType_string = "insTab";
      default : io_inputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_respType)
      LockRespType_grant : io_inputs_1_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_1_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_1_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_1_payload_respType_string = "release_1";
      default : io_inputs_1_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_lkType)
      LkT_rd : io_inputs_2_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_2_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_2_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_2_payload_lkType_string = "insTab";
      default : io_inputs_2_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_respType)
      LockRespType_grant : io_inputs_2_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_2_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_2_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_2_payload_respType_string = "release_1";
      default : io_inputs_2_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_3_payload_lkType)
      LkT_rd : io_inputs_3_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_3_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_3_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_3_payload_lkType_string = "insTab";
      default : io_inputs_3_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_3_payload_respType)
      LockRespType_grant : io_inputs_3_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_3_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_3_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_3_payload_respType_string = "release_1";
      default : io_inputs_3_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_4_payload_lkType)
      LkT_rd : io_inputs_4_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_4_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_4_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_4_payload_lkType_string = "insTab";
      default : io_inputs_4_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_4_payload_respType)
      LockRespType_grant : io_inputs_4_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_4_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_4_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_4_payload_respType_string = "release_1";
      default : io_inputs_4_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_5_payload_lkType)
      LkT_rd : io_inputs_5_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_5_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_5_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_5_payload_lkType_string = "insTab";
      default : io_inputs_5_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_5_payload_respType)
      LockRespType_grant : io_inputs_5_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_5_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_5_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_5_payload_respType_string = "release_1";
      default : io_inputs_5_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_6_payload_lkType)
      LkT_rd : io_inputs_6_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_6_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_6_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_6_payload_lkType_string = "insTab";
      default : io_inputs_6_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_6_payload_respType)
      LockRespType_grant : io_inputs_6_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_6_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_6_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_6_payload_respType_string = "release_1";
      default : io_inputs_6_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_7_payload_lkType)
      LkT_rd : io_inputs_7_payload_lkType_string = "rd    ";
      LkT_wr : io_inputs_7_payload_lkType_string = "wr    ";
      LkT_raw : io_inputs_7_payload_lkType_string = "raw   ";
      LkT_insTab : io_inputs_7_payload_lkType_string = "insTab";
      default : io_inputs_7_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_7_payload_respType)
      LockRespType_grant : io_inputs_7_payload_respType_string = "grant    ";
      LockRespType_abort : io_inputs_7_payload_respType_string = "abort    ";
      LockRespType_waiting : io_inputs_7_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_inputs_7_payload_respType_string = "release_1";
      default : io_inputs_7_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_lkType)
      LkT_rd : io_output_payload_lkType_string = "rd    ";
      LkT_wr : io_output_payload_lkType_string = "wr    ";
      LkT_raw : io_output_payload_lkType_string = "raw   ";
      LkT_insTab : io_output_payload_lkType_string = "insTab";
      default : io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_respType)
      LockRespType_grant : io_output_payload_respType_string = "grant    ";
      LockRespType_abort : io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_output_payload_respType_string = "release_1";
      default : io_output_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_lkType)
      LkT_rd : _zz_io_output_payload_lkType_string = "rd    ";
      LkT_wr : _zz_io_output_payload_lkType_string = "wr    ";
      LkT_raw : _zz_io_output_payload_lkType_string = "raw   ";
      LkT_insTab : _zz_io_output_payload_lkType_string = "insTab";
      default : _zz_io_output_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_respType)
      LockRespType_grant : _zz_io_output_payload_respType_string = "grant    ";
      LockRespType_abort : _zz_io_output_payload_respType_string = "abort    ";
      LockRespType_waiting : _zz_io_output_payload_respType_string = "waiting  ";
      LockRespType_release_1 : _zz_io_output_payload_respType_string = "release_1";
      default : _zz_io_output_payload_respType_string = "?????????";
    endcase
  end
  `endif

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign maskRouted_4 = (locked ? maskLocked_4 : maskProposal_4);
  assign maskRouted_5 = (locked ? maskLocked_5 : maskProposal_5);
  assign maskRouted_6 = (locked ? maskLocked_6 : maskProposal_6);
  assign maskRouted_7 = (locked ? maskLocked_7 : maskProposal_7);
  assign _zz_maskProposal_0 = {io_inputs_7_valid,{io_inputs_6_valid,{io_inputs_5_valid,{io_inputs_4_valid,{io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}}}}}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[15 : 8] | _zz_maskProposal_0_2[7 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign maskProposal_3 = _zz_maskProposal_0_3[3];
  assign maskProposal_4 = _zz_maskProposal_0_3[4];
  assign maskProposal_5 = _zz_maskProposal_0_3[5];
  assign maskProposal_6 = _zz_maskProposal_0_3[6];
  assign maskProposal_7 = _zz_maskProposal_0_3[7];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((((((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3)) || (io_inputs_4_valid && maskRouted_4)) || (io_inputs_5_valid && maskRouted_5)) || (io_inputs_6_valid && maskRouted_6)) || (io_inputs_7_valid && maskRouted_7));
  assign _zz_io_output_payload_nId = (((maskRouted_1 || maskRouted_3) || maskRouted_5) || maskRouted_7);
  assign _zz_io_output_payload_nId_1 = (((maskRouted_2 || maskRouted_3) || maskRouted_6) || maskRouted_7);
  assign _zz_io_output_payload_nId_2 = (((maskRouted_4 || maskRouted_5) || maskRouted_6) || maskRouted_7);
  assign _zz_io_output_payload_nId_3 = {_zz_io_output_payload_nId_2,{_zz_io_output_payload_nId_1,_zz_io_output_payload_nId}};
  assign _zz_io_output_payload_lkType = _zz__zz_io_output_payload_lkType;
  assign _zz_io_output_payload_respType = _zz__zz_io_output_payload_respType;
  assign io_output_payload_nId = _zz_io_output_payload_nId_4;
  assign io_output_payload_tId = _zz_io_output_payload_tId;
  assign io_output_payload_tabId = _zz_io_output_payload_tabId;
  assign io_output_payload_snId = _zz_io_output_payload_snId;
  assign io_output_payload_txnId = _zz_io_output_payload_txnId;
  assign io_output_payload_lkType = _zz_io_output_payload_lkType;
  assign io_output_payload_lkRelease = _zz_io_output_payload_lkRelease;
  assign io_output_payload_txnAbt = _zz_io_output_payload_txnAbt;
  assign io_output_payload_lkIdx = _zz_io_output_payload_lkIdx;
  assign io_output_payload_wLen = _zz_io_output_payload_wLen;
  assign io_output_payload_respType = _zz_io_output_payload_respType;
  assign io_output_payload_lkWaited = _zz_io_output_payload_lkWaited;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_inputs_3_ready = (maskRouted_3 && io_output_ready);
  assign io_inputs_4_ready = (maskRouted_4 && io_output_ready);
  assign io_inputs_5_ready = (maskRouted_5 && io_output_ready);
  assign io_inputs_6_ready = (maskRouted_6 && io_output_ready);
  assign io_inputs_7_ready = (maskRouted_7 && io_output_ready);
  assign io_chosenOH = {maskRouted_7,{maskRouted_6,{maskRouted_5,{maskRouted_4,{maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}}}}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = io_chosenOH[5];
  assign _zz_io_chosen_2 = io_chosenOH[6];
  assign _zz_io_chosen_3 = io_chosenOH[7];
  assign _zz_io_chosen_4 = (((io_chosenOH[1] || _zz_io_chosen) || _zz_io_chosen_1) || _zz_io_chosen_3);
  assign _zz_io_chosen_5 = (((io_chosenOH[2] || _zz_io_chosen) || _zz_io_chosen_2) || _zz_io_chosen_3);
  assign _zz_io_chosen_6 = (((io_chosenOH[4] || _zz_io_chosen_1) || _zz_io_chosen_2) || _zz_io_chosen_3);
  assign io_chosen = {_zz_io_chosen_6,{_zz_io_chosen_5,_zz_io_chosen_4}};
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b0;
      maskLocked_3 <= 1'b0;
      maskLocked_4 <= 1'b0;
      maskLocked_5 <= 1'b0;
      maskLocked_6 <= 1'b0;
      maskLocked_7 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
        maskLocked_3 <= maskRouted_3;
        maskLocked_4 <= maskRouted_4;
        maskLocked_5 <= maskRouted_5;
        maskLocked_6 <= maskRouted_6;
        maskLocked_7 <= maskRouted_7;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamDemux_1 (
  input      [2:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [0:0]    io_input_payload_nId,
  input      [18:0]   io_input_payload_tId,
  input      [2:0]    io_input_payload_tabId,
  input      [0:0]    io_input_payload_snId,
  input      [5:0]    io_input_payload_txnId,
  input      [1:0]    io_input_payload_lkType,
  input               io_input_payload_lkRelease,
  input               io_input_payload_txnTimeOut,
  input               io_input_payload_txnAbt,
  input      [5:0]    io_input_payload_lkIdx,
  input      [2:0]    io_input_payload_wLen,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [0:0]    io_outputs_0_payload_nId,
  output     [18:0]   io_outputs_0_payload_tId,
  output     [2:0]    io_outputs_0_payload_tabId,
  output     [0:0]    io_outputs_0_payload_snId,
  output     [5:0]    io_outputs_0_payload_txnId,
  output     [1:0]    io_outputs_0_payload_lkType,
  output              io_outputs_0_payload_lkRelease,
  output              io_outputs_0_payload_txnTimeOut,
  output              io_outputs_0_payload_txnAbt,
  output     [5:0]    io_outputs_0_payload_lkIdx,
  output     [2:0]    io_outputs_0_payload_wLen,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [0:0]    io_outputs_1_payload_nId,
  output     [18:0]   io_outputs_1_payload_tId,
  output     [2:0]    io_outputs_1_payload_tabId,
  output     [0:0]    io_outputs_1_payload_snId,
  output     [5:0]    io_outputs_1_payload_txnId,
  output     [1:0]    io_outputs_1_payload_lkType,
  output              io_outputs_1_payload_lkRelease,
  output              io_outputs_1_payload_txnTimeOut,
  output              io_outputs_1_payload_txnAbt,
  output     [5:0]    io_outputs_1_payload_lkIdx,
  output     [2:0]    io_outputs_1_payload_wLen,
  output reg          io_outputs_2_valid,
  input               io_outputs_2_ready,
  output     [0:0]    io_outputs_2_payload_nId,
  output     [18:0]   io_outputs_2_payload_tId,
  output     [2:0]    io_outputs_2_payload_tabId,
  output     [0:0]    io_outputs_2_payload_snId,
  output     [5:0]    io_outputs_2_payload_txnId,
  output     [1:0]    io_outputs_2_payload_lkType,
  output              io_outputs_2_payload_lkRelease,
  output              io_outputs_2_payload_txnTimeOut,
  output              io_outputs_2_payload_txnAbt,
  output     [5:0]    io_outputs_2_payload_lkIdx,
  output     [2:0]    io_outputs_2_payload_wLen,
  output reg          io_outputs_3_valid,
  input               io_outputs_3_ready,
  output     [0:0]    io_outputs_3_payload_nId,
  output     [18:0]   io_outputs_3_payload_tId,
  output     [2:0]    io_outputs_3_payload_tabId,
  output     [0:0]    io_outputs_3_payload_snId,
  output     [5:0]    io_outputs_3_payload_txnId,
  output     [1:0]    io_outputs_3_payload_lkType,
  output              io_outputs_3_payload_lkRelease,
  output              io_outputs_3_payload_txnTimeOut,
  output              io_outputs_3_payload_txnAbt,
  output     [5:0]    io_outputs_3_payload_lkIdx,
  output     [2:0]    io_outputs_3_payload_wLen,
  output reg          io_outputs_4_valid,
  input               io_outputs_4_ready,
  output     [0:0]    io_outputs_4_payload_nId,
  output     [18:0]   io_outputs_4_payload_tId,
  output     [2:0]    io_outputs_4_payload_tabId,
  output     [0:0]    io_outputs_4_payload_snId,
  output     [5:0]    io_outputs_4_payload_txnId,
  output     [1:0]    io_outputs_4_payload_lkType,
  output              io_outputs_4_payload_lkRelease,
  output              io_outputs_4_payload_txnTimeOut,
  output              io_outputs_4_payload_txnAbt,
  output     [5:0]    io_outputs_4_payload_lkIdx,
  output     [2:0]    io_outputs_4_payload_wLen,
  output reg          io_outputs_5_valid,
  input               io_outputs_5_ready,
  output     [0:0]    io_outputs_5_payload_nId,
  output     [18:0]   io_outputs_5_payload_tId,
  output     [2:0]    io_outputs_5_payload_tabId,
  output     [0:0]    io_outputs_5_payload_snId,
  output     [5:0]    io_outputs_5_payload_txnId,
  output     [1:0]    io_outputs_5_payload_lkType,
  output              io_outputs_5_payload_lkRelease,
  output              io_outputs_5_payload_txnTimeOut,
  output              io_outputs_5_payload_txnAbt,
  output     [5:0]    io_outputs_5_payload_lkIdx,
  output     [2:0]    io_outputs_5_payload_wLen,
  output reg          io_outputs_6_valid,
  input               io_outputs_6_ready,
  output     [0:0]    io_outputs_6_payload_nId,
  output     [18:0]   io_outputs_6_payload_tId,
  output     [2:0]    io_outputs_6_payload_tabId,
  output     [0:0]    io_outputs_6_payload_snId,
  output     [5:0]    io_outputs_6_payload_txnId,
  output     [1:0]    io_outputs_6_payload_lkType,
  output              io_outputs_6_payload_lkRelease,
  output              io_outputs_6_payload_txnTimeOut,
  output              io_outputs_6_payload_txnAbt,
  output     [5:0]    io_outputs_6_payload_lkIdx,
  output     [2:0]    io_outputs_6_payload_wLen,
  output reg          io_outputs_7_valid,
  input               io_outputs_7_ready,
  output     [0:0]    io_outputs_7_payload_nId,
  output     [18:0]   io_outputs_7_payload_tId,
  output     [2:0]    io_outputs_7_payload_tabId,
  output     [0:0]    io_outputs_7_payload_snId,
  output     [5:0]    io_outputs_7_payload_txnId,
  output     [1:0]    io_outputs_7_payload_lkType,
  output              io_outputs_7_payload_lkRelease,
  output              io_outputs_7_payload_txnTimeOut,
  output              io_outputs_7_payload_txnAbt,
  output     [5:0]    io_outputs_7_payload_lkIdx,
  output     [2:0]    io_outputs_7_payload_wLen
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire                when_Stream_l881;
  wire                when_Stream_l881_1;
  wire                when_Stream_l881_2;
  wire                when_Stream_l881_3;
  wire                when_Stream_l881_4;
  wire                when_Stream_l881_5;
  wire                when_Stream_l881_6;
  wire                when_Stream_l881_7;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_lkType_string;
  reg [47:0] io_outputs_0_payload_lkType_string;
  reg [47:0] io_outputs_1_payload_lkType_string;
  reg [47:0] io_outputs_2_payload_lkType_string;
  reg [47:0] io_outputs_3_payload_lkType_string;
  reg [47:0] io_outputs_4_payload_lkType_string;
  reg [47:0] io_outputs_5_payload_lkType_string;
  reg [47:0] io_outputs_6_payload_lkType_string;
  reg [47:0] io_outputs_7_payload_lkType_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_lkType)
      LkT_rd : io_input_payload_lkType_string = "rd    ";
      LkT_wr : io_input_payload_lkType_string = "wr    ";
      LkT_raw : io_input_payload_lkType_string = "raw   ";
      LkT_insTab : io_input_payload_lkType_string = "insTab";
      default : io_input_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_lkType)
      LkT_rd : io_outputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_0_payload_lkType_string = "insTab";
      default : io_outputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_lkType)
      LkT_rd : io_outputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_1_payload_lkType_string = "insTab";
      default : io_outputs_1_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_2_payload_lkType)
      LkT_rd : io_outputs_2_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_2_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_2_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_2_payload_lkType_string = "insTab";
      default : io_outputs_2_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_3_payload_lkType)
      LkT_rd : io_outputs_3_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_3_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_3_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_3_payload_lkType_string = "insTab";
      default : io_outputs_3_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_4_payload_lkType)
      LkT_rd : io_outputs_4_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_4_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_4_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_4_payload_lkType_string = "insTab";
      default : io_outputs_4_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_5_payload_lkType)
      LkT_rd : io_outputs_5_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_5_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_5_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_5_payload_lkType_string = "insTab";
      default : io_outputs_5_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_6_payload_lkType)
      LkT_rd : io_outputs_6_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_6_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_6_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_6_payload_lkType_string = "insTab";
      default : io_outputs_6_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_7_payload_lkType)
      LkT_rd : io_outputs_7_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_7_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_7_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_7_payload_lkType_string = "insTab";
      default : io_outputs_7_payload_lkType_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l881) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l881_1) begin
      io_input_ready = io_outputs_1_ready;
    end
    if(!when_Stream_l881_2) begin
      io_input_ready = io_outputs_2_ready;
    end
    if(!when_Stream_l881_3) begin
      io_input_ready = io_outputs_3_ready;
    end
    if(!when_Stream_l881_4) begin
      io_input_ready = io_outputs_4_ready;
    end
    if(!when_Stream_l881_5) begin
      io_input_ready = io_outputs_5_ready;
    end
    if(!when_Stream_l881_6) begin
      io_input_ready = io_outputs_6_ready;
    end
    if(!when_Stream_l881_7) begin
      io_input_ready = io_outputs_7_ready;
    end
  end

  assign io_outputs_0_payload_nId = io_input_payload_nId;
  assign io_outputs_0_payload_tId = io_input_payload_tId;
  assign io_outputs_0_payload_tabId = io_input_payload_tabId;
  assign io_outputs_0_payload_snId = io_input_payload_snId;
  assign io_outputs_0_payload_txnId = io_input_payload_txnId;
  assign io_outputs_0_payload_lkType = io_input_payload_lkType;
  assign io_outputs_0_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_0_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_0_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_0_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_0_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881 = (3'b000 != io_select);
  always @(*) begin
    if(when_Stream_l881) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_nId = io_input_payload_nId;
  assign io_outputs_1_payload_tId = io_input_payload_tId;
  assign io_outputs_1_payload_tabId = io_input_payload_tabId;
  assign io_outputs_1_payload_snId = io_input_payload_snId;
  assign io_outputs_1_payload_txnId = io_input_payload_txnId;
  assign io_outputs_1_payload_lkType = io_input_payload_lkType;
  assign io_outputs_1_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_1_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_1_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_1_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_1_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_1 = (3'b001 != io_select);
  always @(*) begin
    if(when_Stream_l881_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end

  assign io_outputs_2_payload_nId = io_input_payload_nId;
  assign io_outputs_2_payload_tId = io_input_payload_tId;
  assign io_outputs_2_payload_tabId = io_input_payload_tabId;
  assign io_outputs_2_payload_snId = io_input_payload_snId;
  assign io_outputs_2_payload_txnId = io_input_payload_txnId;
  assign io_outputs_2_payload_lkType = io_input_payload_lkType;
  assign io_outputs_2_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_2_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_2_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_2_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_2_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_2 = (3'b010 != io_select);
  always @(*) begin
    if(when_Stream_l881_2) begin
      io_outputs_2_valid = 1'b0;
    end else begin
      io_outputs_2_valid = io_input_valid;
    end
  end

  assign io_outputs_3_payload_nId = io_input_payload_nId;
  assign io_outputs_3_payload_tId = io_input_payload_tId;
  assign io_outputs_3_payload_tabId = io_input_payload_tabId;
  assign io_outputs_3_payload_snId = io_input_payload_snId;
  assign io_outputs_3_payload_txnId = io_input_payload_txnId;
  assign io_outputs_3_payload_lkType = io_input_payload_lkType;
  assign io_outputs_3_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_3_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_3_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_3_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_3_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_3 = (3'b011 != io_select);
  always @(*) begin
    if(when_Stream_l881_3) begin
      io_outputs_3_valid = 1'b0;
    end else begin
      io_outputs_3_valid = io_input_valid;
    end
  end

  assign io_outputs_4_payload_nId = io_input_payload_nId;
  assign io_outputs_4_payload_tId = io_input_payload_tId;
  assign io_outputs_4_payload_tabId = io_input_payload_tabId;
  assign io_outputs_4_payload_snId = io_input_payload_snId;
  assign io_outputs_4_payload_txnId = io_input_payload_txnId;
  assign io_outputs_4_payload_lkType = io_input_payload_lkType;
  assign io_outputs_4_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_4_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_4_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_4_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_4_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_4 = (3'b100 != io_select);
  always @(*) begin
    if(when_Stream_l881_4) begin
      io_outputs_4_valid = 1'b0;
    end else begin
      io_outputs_4_valid = io_input_valid;
    end
  end

  assign io_outputs_5_payload_nId = io_input_payload_nId;
  assign io_outputs_5_payload_tId = io_input_payload_tId;
  assign io_outputs_5_payload_tabId = io_input_payload_tabId;
  assign io_outputs_5_payload_snId = io_input_payload_snId;
  assign io_outputs_5_payload_txnId = io_input_payload_txnId;
  assign io_outputs_5_payload_lkType = io_input_payload_lkType;
  assign io_outputs_5_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_5_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_5_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_5_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_5_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_5 = (3'b101 != io_select);
  always @(*) begin
    if(when_Stream_l881_5) begin
      io_outputs_5_valid = 1'b0;
    end else begin
      io_outputs_5_valid = io_input_valid;
    end
  end

  assign io_outputs_6_payload_nId = io_input_payload_nId;
  assign io_outputs_6_payload_tId = io_input_payload_tId;
  assign io_outputs_6_payload_tabId = io_input_payload_tabId;
  assign io_outputs_6_payload_snId = io_input_payload_snId;
  assign io_outputs_6_payload_txnId = io_input_payload_txnId;
  assign io_outputs_6_payload_lkType = io_input_payload_lkType;
  assign io_outputs_6_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_6_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_6_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_6_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_6_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_6 = (3'b110 != io_select);
  always @(*) begin
    if(when_Stream_l881_6) begin
      io_outputs_6_valid = 1'b0;
    end else begin
      io_outputs_6_valid = io_input_valid;
    end
  end

  assign io_outputs_7_payload_nId = io_input_payload_nId;
  assign io_outputs_7_payload_tId = io_input_payload_tId;
  assign io_outputs_7_payload_tabId = io_input_payload_tabId;
  assign io_outputs_7_payload_snId = io_input_payload_snId;
  assign io_outputs_7_payload_txnId = io_input_payload_txnId;
  assign io_outputs_7_payload_lkType = io_input_payload_lkType;
  assign io_outputs_7_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_7_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_7_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_7_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_7_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_7 = (3'b111 != io_select);
  always @(*) begin
    if(when_Stream_l881_7) begin
      io_outputs_7_valid = 1'b0;
    end else begin
      io_outputs_7_valid = io_input_valid;
    end
  end


endmodule

module StreamDemux (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [0:0]    io_input_payload_nId,
  input      [21:0]   io_input_payload_tId,
  input      [2:0]    io_input_payload_tabId,
  input      [0:0]    io_input_payload_snId,
  input      [5:0]    io_input_payload_txnId,
  input      [1:0]    io_input_payload_lkType,
  input               io_input_payload_lkRelease,
  input               io_input_payload_txnTimeOut,
  input               io_input_payload_txnAbt,
  input      [5:0]    io_input_payload_lkIdx,
  input      [2:0]    io_input_payload_wLen,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [0:0]    io_outputs_0_payload_nId,
  output     [21:0]   io_outputs_0_payload_tId,
  output     [2:0]    io_outputs_0_payload_tabId,
  output     [0:0]    io_outputs_0_payload_snId,
  output     [5:0]    io_outputs_0_payload_txnId,
  output     [1:0]    io_outputs_0_payload_lkType,
  output              io_outputs_0_payload_lkRelease,
  output              io_outputs_0_payload_txnTimeOut,
  output              io_outputs_0_payload_txnAbt,
  output     [5:0]    io_outputs_0_payload_lkIdx,
  output     [2:0]    io_outputs_0_payload_wLen,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [0:0]    io_outputs_1_payload_nId,
  output     [21:0]   io_outputs_1_payload_tId,
  output     [2:0]    io_outputs_1_payload_tabId,
  output     [0:0]    io_outputs_1_payload_snId,
  output     [5:0]    io_outputs_1_payload_txnId,
  output     [1:0]    io_outputs_1_payload_lkType,
  output              io_outputs_1_payload_lkRelease,
  output              io_outputs_1_payload_txnTimeOut,
  output              io_outputs_1_payload_txnAbt,
  output     [5:0]    io_outputs_1_payload_lkIdx,
  output     [2:0]    io_outputs_1_payload_wLen
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;

  wire                when_Stream_l881;
  wire                when_Stream_l881_1;
  `ifndef SYNTHESIS
  reg [47:0] io_input_payload_lkType_string;
  reg [47:0] io_outputs_0_payload_lkType_string;
  reg [47:0] io_outputs_1_payload_lkType_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_lkType)
      LkT_rd : io_input_payload_lkType_string = "rd    ";
      LkT_wr : io_input_payload_lkType_string = "wr    ";
      LkT_raw : io_input_payload_lkType_string = "raw   ";
      LkT_insTab : io_input_payload_lkType_string = "insTab";
      default : io_input_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_lkType)
      LkT_rd : io_outputs_0_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_0_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_0_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_0_payload_lkType_string = "insTab";
      default : io_outputs_0_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_lkType)
      LkT_rd : io_outputs_1_payload_lkType_string = "rd    ";
      LkT_wr : io_outputs_1_payload_lkType_string = "wr    ";
      LkT_raw : io_outputs_1_payload_lkType_string = "raw   ";
      LkT_insTab : io_outputs_1_payload_lkType_string = "insTab";
      default : io_outputs_1_payload_lkType_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l881) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l881_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_nId = io_input_payload_nId;
  assign io_outputs_0_payload_tId = io_input_payload_tId;
  assign io_outputs_0_payload_tabId = io_input_payload_tabId;
  assign io_outputs_0_payload_snId = io_input_payload_snId;
  assign io_outputs_0_payload_txnId = io_input_payload_txnId;
  assign io_outputs_0_payload_lkType = io_input_payload_lkType;
  assign io_outputs_0_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_0_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_0_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_0_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_0_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l881) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_nId = io_input_payload_nId;
  assign io_outputs_1_payload_tId = io_input_payload_tId;
  assign io_outputs_1_payload_tabId = io_input_payload_tabId;
  assign io_outputs_1_payload_snId = io_input_payload_snId;
  assign io_outputs_1_payload_txnId = io_input_payload_txnId;
  assign io_outputs_1_payload_lkType = io_input_payload_lkType;
  assign io_outputs_1_payload_lkRelease = io_input_payload_lkRelease;
  assign io_outputs_1_payload_txnTimeOut = io_input_payload_txnTimeOut;
  assign io_outputs_1_payload_txnAbt = io_input_payload_txnAbt;
  assign io_outputs_1_payload_lkIdx = io_input_payload_lkIdx;
  assign io_outputs_1_payload_wLen = io_input_payload_wLen;
  assign when_Stream_l881_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l881_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module LockTableBW_7 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_7_BOOT = 4'd0;
  localparam htFsm_enumDef_7_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_7_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_7_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_7_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_7_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_7_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_7_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_7_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_7_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_7_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_7_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_7_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_7_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_7_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_7_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_7_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_7_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_7_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_7_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_7_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_7_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_7_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_7_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_7_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_7_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_7_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_7_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_7_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_7_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_7_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_7_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_7_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_7_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_7_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_7_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_7_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_7_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_7_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
      end
      htFsm_enumDef_7_HTINSRESP : begin
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_7_LKRESP) || (htFsm_stateReg == htFsm_enumDef_7_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_7_HTINSRESP;
        end
      end
      htFsm_enumDef_7_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_7_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_7_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_7_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_7_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_7_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_7_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_7_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_7_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_7_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_7_HTDELRESP;
        end
      end
      htFsm_enumDef_7_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_7_LKRESP;
        end
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_7_LLPUSHRESP;
        end
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_7_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_7_LKRESP;
          end
        end
      end
      htFsm_enumDef_7_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_7_LLPOPRESP;
        end
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_7_LKRESP;
        end
      end
      htFsm_enumDef_7_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_7_LLDELRESP;
        end
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_7_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_7_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_7_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_7_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_7_LLPOPCMD;
        end
      end
      htFsm_enumDef_7_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_7_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_7_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_7_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_7_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_7_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_7_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_7_HTDELCMD : begin
      end
      htFsm_enumDef_7_HTDELRESP : begin
      end
      htFsm_enumDef_7_LLPUSHCMD : begin
      end
      htFsm_enumDef_7_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_7_LLPOPCMD : begin
      end
      htFsm_enumDef_7_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_7_LLDELCMD : begin
      end
      htFsm_enumDef_7_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_7_LKRESPPOP : begin
      end
      htFsm_enumDef_7_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_7_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_6 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_6_BOOT = 4'd0;
  localparam htFsm_enumDef_6_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_6_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_6_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_6_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_6_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_6_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_6_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_6_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_6_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_6_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_6_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_6_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_6_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_6_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_6_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_6_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_6_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_6_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_6_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_6_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_6_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_6_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_6_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_6_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_6_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_6_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_6_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_6_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_6_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_6_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_6_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_6_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_6_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_6_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_6_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_6_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_6_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_6_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
      end
      htFsm_enumDef_6_HTINSRESP : begin
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_6_LKRESP) || (htFsm_stateReg == htFsm_enumDef_6_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_6_HTINSRESP;
        end
      end
      htFsm_enumDef_6_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_6_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_6_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_6_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_6_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_6_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_6_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_6_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_6_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_6_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_6_HTDELRESP;
        end
      end
      htFsm_enumDef_6_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_6_LKRESP;
        end
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_6_LLPUSHRESP;
        end
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_6_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_6_LKRESP;
          end
        end
      end
      htFsm_enumDef_6_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_6_LLPOPRESP;
        end
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_6_LKRESP;
        end
      end
      htFsm_enumDef_6_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_6_LLDELRESP;
        end
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_6_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_6_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_6_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_6_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_6_LLPOPCMD;
        end
      end
      htFsm_enumDef_6_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_6_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_6_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_6_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_6_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_6_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_6_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_6_HTDELCMD : begin
      end
      htFsm_enumDef_6_HTDELRESP : begin
      end
      htFsm_enumDef_6_LLPUSHCMD : begin
      end
      htFsm_enumDef_6_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_6_LLPOPCMD : begin
      end
      htFsm_enumDef_6_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_6_LLDELCMD : begin
      end
      htFsm_enumDef_6_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_6_LKRESPPOP : begin
      end
      htFsm_enumDef_6_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_6_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_5 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_5_BOOT = 4'd0;
  localparam htFsm_enumDef_5_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_5_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_5_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_5_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_5_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_5_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_5_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_5_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_5_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_5_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_5_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_5_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_5_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_5_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_5_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_5_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_5_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_5_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_5_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_5_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_5_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_5_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_5_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_5_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_5_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_5_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_5_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_5_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_5_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_5_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_5_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_5_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_5_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_5_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_5_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_5_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_5_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_5_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
      end
      htFsm_enumDef_5_HTINSRESP : begin
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_5_LKRESP) || (htFsm_stateReg == htFsm_enumDef_5_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_5_HTINSRESP;
        end
      end
      htFsm_enumDef_5_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_5_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_5_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_5_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_5_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_5_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_5_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_5_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_5_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_5_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_5_HTDELRESP;
        end
      end
      htFsm_enumDef_5_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_5_LKRESP;
        end
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_5_LLPUSHRESP;
        end
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_5_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_5_LKRESP;
          end
        end
      end
      htFsm_enumDef_5_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_5_LLPOPRESP;
        end
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_5_LKRESP;
        end
      end
      htFsm_enumDef_5_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_5_LLDELRESP;
        end
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_5_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_5_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_5_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_5_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_5_LLPOPCMD;
        end
      end
      htFsm_enumDef_5_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_5_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_5_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_5_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_5_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_5_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_5_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_5_HTDELCMD : begin
      end
      htFsm_enumDef_5_HTDELRESP : begin
      end
      htFsm_enumDef_5_LLPUSHCMD : begin
      end
      htFsm_enumDef_5_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_5_LLPOPCMD : begin
      end
      htFsm_enumDef_5_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_5_LLDELCMD : begin
      end
      htFsm_enumDef_5_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_5_LKRESPPOP : begin
      end
      htFsm_enumDef_5_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_5_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_4 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_4_BOOT = 4'd0;
  localparam htFsm_enumDef_4_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_4_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_4_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_4_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_4_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_4_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_4_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_4_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_4_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_4_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_4_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_4_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_4_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_4_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_4_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_4_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_4_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_4_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_4_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_4_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_4_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_4_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_4_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_4_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_4_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_4_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_4_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_4_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_4_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_4_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_4_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_4_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_4_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_4_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_4_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_4_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_4_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_4_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
      end
      htFsm_enumDef_4_HTINSRESP : begin
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_4_LKRESP) || (htFsm_stateReg == htFsm_enumDef_4_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_4_HTINSRESP;
        end
      end
      htFsm_enumDef_4_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_4_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_4_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_4_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_4_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_4_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_4_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_4_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_4_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_4_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_4_HTDELRESP;
        end
      end
      htFsm_enumDef_4_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_4_LKRESP;
        end
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_4_LLPUSHRESP;
        end
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_4_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_4_LKRESP;
          end
        end
      end
      htFsm_enumDef_4_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_4_LLPOPRESP;
        end
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_4_LKRESP;
        end
      end
      htFsm_enumDef_4_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_4_LLDELRESP;
        end
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_4_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_4_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_4_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_4_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_4_LLPOPCMD;
        end
      end
      htFsm_enumDef_4_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_4_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_4_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_4_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_4_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_4_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_4_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_4_HTDELCMD : begin
      end
      htFsm_enumDef_4_HTDELRESP : begin
      end
      htFsm_enumDef_4_LLPUSHCMD : begin
      end
      htFsm_enumDef_4_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_4_LLPOPCMD : begin
      end
      htFsm_enumDef_4_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_4_LLDELCMD : begin
      end
      htFsm_enumDef_4_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_4_LKRESPPOP : begin
      end
      htFsm_enumDef_4_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_4_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_3 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_3_BOOT = 4'd0;
  localparam htFsm_enumDef_3_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_3_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_3_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_3_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_3_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_3_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_3_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_3_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_3_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_3_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_3_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_3_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_3_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_3_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_3_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_3_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_3_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_3_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_3_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_3_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_3_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_3_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_3_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_3_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_3_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_3_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_3_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_3_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_3_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_3_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_3_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_3_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_3_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_3_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_3_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_3_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_3_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_3_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
      end
      htFsm_enumDef_3_HTINSRESP : begin
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_3_LKRESP) || (htFsm_stateReg == htFsm_enumDef_3_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_3_HTINSRESP;
        end
      end
      htFsm_enumDef_3_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_3_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_3_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_3_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_3_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_3_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_3_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_3_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_3_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_3_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_3_HTDELRESP;
        end
      end
      htFsm_enumDef_3_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_3_LKRESP;
        end
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_3_LLPUSHRESP;
        end
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_3_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_3_LKRESP;
          end
        end
      end
      htFsm_enumDef_3_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_3_LLPOPRESP;
        end
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_3_LKRESP;
        end
      end
      htFsm_enumDef_3_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_3_LLDELRESP;
        end
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_3_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_3_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_3_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_3_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_3_LLPOPCMD;
        end
      end
      htFsm_enumDef_3_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_3_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_3_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_3_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_3_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_3_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_3_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_3_HTDELCMD : begin
      end
      htFsm_enumDef_3_HTDELRESP : begin
      end
      htFsm_enumDef_3_LLPUSHCMD : begin
      end
      htFsm_enumDef_3_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_3_LLPOPCMD : begin
      end
      htFsm_enumDef_3_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_3_LLDELCMD : begin
      end
      htFsm_enumDef_3_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_3_LKRESPPOP : begin
      end
      htFsm_enumDef_3_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_3_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_2 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_2_BOOT = 4'd0;
  localparam htFsm_enumDef_2_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_2_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_2_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_2_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_2_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_2_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_2_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_2_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_2_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_2_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_2_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_2_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_2_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_2_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_2_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_2_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_2_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_2_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_2_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_2_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_2_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_2_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_2_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_2_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_2_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_2_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_2_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_2_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_2_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_2_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_2_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_2_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_2_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_2_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_2_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_2_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_2_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_2_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
      end
      htFsm_enumDef_2_HTINSRESP : begin
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_2_LKRESP) || (htFsm_stateReg == htFsm_enumDef_2_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_2_HTINSRESP;
        end
      end
      htFsm_enumDef_2_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_2_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_2_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_2_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_2_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_2_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_2_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_2_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_2_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_2_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_2_HTDELRESP;
        end
      end
      htFsm_enumDef_2_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_2_LKRESP;
        end
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_2_LLPUSHRESP;
        end
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_2_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_2_LKRESP;
          end
        end
      end
      htFsm_enumDef_2_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_2_LLPOPRESP;
        end
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_2_LKRESP;
        end
      end
      htFsm_enumDef_2_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_2_LLDELRESP;
        end
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_2_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_2_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_2_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_2_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_2_LLPOPCMD;
        end
      end
      htFsm_enumDef_2_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_2_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_2_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_2_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_2_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_2_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_2_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_2_HTDELCMD : begin
      end
      htFsm_enumDef_2_HTDELRESP : begin
      end
      htFsm_enumDef_2_LLPUSHCMD : begin
      end
      htFsm_enumDef_2_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_2_LLPOPCMD : begin
      end
      htFsm_enumDef_2_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_2_LLDELCMD : begin
      end
      htFsm_enumDef_2_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_2_LKRESPPOP : begin
      end
      htFsm_enumDef_2_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_2_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW_1 (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_1_BOOT = 4'd0;
  localparam htFsm_enumDef_1_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_1_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_1_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_1_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_1_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_1_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_1_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_1_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_1_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_1_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_1_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_1_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_1_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_1_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_1_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_1_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_1_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_1_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_1_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_1_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_1_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_1_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_1_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_1_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_1_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_1_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_1_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_1_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_1_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_1_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_1_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_1_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_1_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_1_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_1_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_1_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_1_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_1_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
      end
      htFsm_enumDef_1_HTINSRESP : begin
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_1_LKRESP) || (htFsm_stateReg == htFsm_enumDef_1_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_1_HTINSRESP;
        end
      end
      htFsm_enumDef_1_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_1_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_1_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_1_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_1_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_1_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_1_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_1_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_1_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_1_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_1_HTDELRESP;
        end
      end
      htFsm_enumDef_1_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_1_LKRESP;
        end
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_1_LLPUSHRESP;
        end
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_1_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_1_LKRESP;
          end
        end
      end
      htFsm_enumDef_1_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_1_LLPOPRESP;
        end
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_1_LKRESP;
        end
      end
      htFsm_enumDef_1_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_1_LLDELRESP;
        end
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_1_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_1_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_1_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_1_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_1_LLPOPCMD;
        end
      end
      htFsm_enumDef_1_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_1_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_1_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_1_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_1_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_1_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_1_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_1_HTDELCMD : begin
      end
      htFsm_enumDef_1_HTDELRESP : begin
      end
      htFsm_enumDef_1_LLPUSHCMD : begin
      end
      htFsm_enumDef_1_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_1_LLPOPCMD : begin
      end
      htFsm_enumDef_1_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_1_LLDELCMD : begin
      end
      htFsm_enumDef_1_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_1_LKRESPPOP : begin
      end
      htFsm_enumDef_1_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_1_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

module LockTableBW (
  input               io_lkReq_valid,
  output reg          io_lkReq_ready,
  input      [0:0]    io_lkReq_payload_nId,
  input      [18:0]   io_lkReq_payload_tId,
  input      [2:0]    io_lkReq_payload_tabId,
  input      [0:0]    io_lkReq_payload_snId,
  input      [5:0]    io_lkReq_payload_txnId,
  input      [1:0]    io_lkReq_payload_lkType,
  input               io_lkReq_payload_lkRelease,
  input               io_lkReq_payload_txnTimeOut,
  input               io_lkReq_payload_txnAbt,
  input      [5:0]    io_lkReq_payload_lkIdx,
  input      [2:0]    io_lkReq_payload_wLen,
  output              io_lkResp_valid,
  input               io_lkResp_ready,
  output     [0:0]    io_lkResp_payload_nId,
  output     [18:0]   io_lkResp_payload_tId,
  output     [2:0]    io_lkResp_payload_tabId,
  output     [0:0]    io_lkResp_payload_snId,
  output     [5:0]    io_lkResp_payload_txnId,
  output     [1:0]    io_lkResp_payload_lkType,
  output              io_lkResp_payload_lkRelease,
  output              io_lkResp_payload_txnAbt,
  output     [5:0]    io_lkResp_payload_lkIdx,
  output     [2:0]    io_lkResp_payload_wLen,
  output     [1:0]    io_lkResp_payload_respType,
  output              io_lkResp_payload_lkWaited,
  input               resetn,
  input               clk
);
  localparam LkT_rd = 2'd0;
  localparam LkT_wr = 2'd1;
  localparam LkT_raw = 2'd2;
  localparam LkT_insTab = 2'd3;
  localparam LockRespType_grant = 2'd0;
  localparam LockRespType_abort = 2'd1;
  localparam LockRespType_waiting = 2'd2;
  localparam LockRespType_release_1 = 2'd3;
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam htFsm_enumDef_BOOT = 4'd0;
  localparam htFsm_enumDef_HTINSCMD = 4'd1;
  localparam htFsm_enumDef_HTINSRESP = 4'd2;
  localparam htFsm_enumDef_HTDELCMD = 4'd3;
  localparam htFsm_enumDef_HTDELRESP = 4'd4;
  localparam htFsm_enumDef_LLPUSHCMD = 4'd5;
  localparam htFsm_enumDef_LLPUSHRESP = 4'd6;
  localparam htFsm_enumDef_LLPOPCMD = 4'd7;
  localparam htFsm_enumDef_LLPOPRESP = 4'd8;
  localparam htFsm_enumDef_LLDELCMD = 4'd9;
  localparam htFsm_enumDef_LLDELRESP = 4'd10;
  localparam htFsm_enumDef_LKRESPPOP = 4'd11;
  localparam htFsm_enumDef_LKRESP = 4'd12;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ht_io_clk_i;
  wire                ht_io_rst_i;
  reg                 ht_io_ht_cmd_if_valid;
  reg        [18:0]   ht_io_ht_cmd_if_payload_key;
  reg        [18:0]   ht_io_ht_cmd_if_payload_value;
  reg        [1:0]    ht_io_ht_cmd_if_payload_opcode;
  reg                 ht_io_update_en;
  reg        [47:0]   ht_io_update_data;
  reg        [8:0]    ht_io_update_addr;
  wire                ll_io_clk_i;
  wire                ll_io_rst_i;
  reg                 ll_io_ll_cmd_if_valid;
  reg        [43:0]   ll_io_ll_cmd_if_payload_key;
  reg        [1:0]    ll_io_ll_cmd_if_payload_opcode;
  reg        [8:0]    ll_io_ll_cmd_if_payload_head_ptr;
  reg                 ll_io_ll_cmd_if_payload_head_ptr_val;
  wire                ht_io_ht_cmd_if_ready;
  wire                ht_io_ht_res_if_valid;
  wire       [47:0]   ht_io_ht_res_if_payload_ram_data;
  wire       [8:0]    ht_io_ht_res_if_payload_find_addr;
  wire       [2:0]    ht_io_ht_res_if_payload_chain_state;
  wire       [18:0]   ht_io_ht_res_if_payload_found_value;
  wire       [7:0]    ht_io_ht_res_if_payload_bucket;
  wire       [2:0]    ht_io_ht_res_if_payload_rescode;
  wire       [1:0]    ht_io_ht_res_if_payload_opcode;
  wire       [18:0]   ht_io_ht_res_if_payload_value;
  wire       [18:0]   ht_io_ht_res_if_payload_key;
  wire                ht_io_ht_clear_ram_done;
  wire                ht_io_dt_clear_ram_done;
  wire                ll_io_ll_cmd_if_ready;
  wire                ll_io_ll_res_if_valid;
  wire       [43:0]   ll_io_ll_res_if_payload_key;
  wire       [1:0]    ll_io_ll_res_if_payload_opcode;
  wire       [2:0]    ll_io_ll_res_if_payload_rescode;
  wire       [2:0]    ll_io_ll_res_if_payload_chain_state;
  wire       [8:0]    ll_io_head_table_if_wr_data_ptr;
  wire                ll_io_head_table_if_wr_data_ptr_val;
  wire                ll_io_head_table_if_wr_en;
  wire                ll_io_clear_ram_done_o;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt;
  wire       [7:0]    _zz_htFsm_htNewRamEntry_ownerCnt_1;
  wire                htFsm_wantExit;
  reg                 htFsm_wantStart;
  wire                htFsm_wantKill;
  reg        [0:0]    htFsm_rLkReq_nId;
  reg        [18:0]   htFsm_rLkReq_tId;
  reg        [2:0]    htFsm_rLkReq_tabId;
  reg        [0:0]    htFsm_rLkReq_snId;
  reg        [5:0]    htFsm_rLkReq_txnId;
  reg        [1:0]    htFsm_rLkReq_lkType;
  reg                 htFsm_rLkReq_lkRelease;
  reg                 htFsm_rLkReq_txnTimeOut;
  reg                 htFsm_rLkReq_txnAbt;
  reg        [5:0]    htFsm_rLkReq_lkIdx;
  reg        [2:0]    htFsm_rLkReq_wLen;
  wire                htFsm_htLkEntry_lkMode;
  wire       [7:0]    htFsm_htLkEntry_ownerCnt;
  wire       [8:0]    htFsm_htLkEntry_waitQPtr;
  wire                htFsm_htLkEntry_waitQPtrVld;
  wire       [18:0]   _zz_htFsm_htLkEntry_lkMode;
  wire                htFsm_htRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htRamEntry_nextPtr;
  wire                htFsm_htRamEntry_lkMode;
  wire       [7:0]    htFsm_htRamEntry_ownerCnt;
  wire       [8:0]    htFsm_htRamEntry_waitQPtr;
  wire                htFsm_htRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htRamEntry_key;
  wire                htFsm_htNewRamEntry_nextPtrVld;
  wire       [8:0]    htFsm_htNewRamEntry_nextPtr;
  reg                 htFsm_htNewRamEntry_lkMode;
  reg        [7:0]    htFsm_htNewRamEntry_ownerCnt;
  reg        [8:0]    htFsm_htNewRamEntry_waitQPtr;
  reg                 htFsm_htNewRamEntry_waitQPtrVld;
  wire       [18:0]   htFsm_htNewRamEntry_key;
  wire       [47:0]   _zz_htFsm_htRamEntry_nextPtrVld;
  wire                ht_io_ht_res_if_fire;
  reg                 htFsm_rHtRamEntry_nextPtrVld;
  reg        [8:0]    htFsm_rHtRamEntry_nextPtr;
  reg                 htFsm_rHtRamEntry_lkMode;
  reg        [7:0]    htFsm_rHtRamEntry_ownerCnt;
  reg        [8:0]    htFsm_rHtRamEntry_waitQPtr;
  reg                 htFsm_rHtRamEntry_waitQPtrVld;
  reg        [18:0]   htFsm_rHtRamEntry_key;
  wire                ht_io_ht_res_if_fire_1;
  reg        [8:0]    htFsm_rHtRamAddr;
  wire                _zz_htFsm_htNewRamEntry_nextPtrVld;
  reg        [1:0]    htFsm_rLkResp;
  reg                 htFsm_rLkWaited;
  wire                htFsm_tryLkEntry_lkMode;
  wire       [7:0]    htFsm_tryLkEntry_ownerCnt;
  wire       [8:0]    htFsm_tryLkEntry_waitQPtr;
  wire                htFsm_tryLkEntry_waitQPtrVld;
  reg        [3:0]    htFsm_stateReg;
  reg        [3:0]    htFsm_stateNext;
  wire                io_lkReq_fire;
  wire                ht_io_ht_res_if_fire_2;
  wire                when_LockTableBW_l109;
  wire                when_LockTableBW_l140;
  wire                ht_io_ht_cmd_if_fire;
  wire                ht_io_ht_res_if_fire_3;
  wire                ll_io_ll_cmd_if_fire;
  wire                ll_io_ll_res_if_fire;
  wire                when_LockTableBW_l184;
  wire                ll_io_ll_cmd_if_fire_1;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType;
  wire       [43:0]   _zz_htFsm_rLkReq_nId;
  wire       [1:0]    _zz_htFsm_rLkReq_lkType_1;
  wire                ll_io_ll_res_if_fire_1;
  wire       [1:0]    _zz_io_ll_cmd_if_payload_key;
  reg                 _zz_io_ll_cmd_if_payload_key_1;
  reg                 _zz_io_ll_cmd_if_payload_key_2;
  reg                 _zz_io_ll_cmd_if_payload_key_3;
  wire                ll_io_ll_cmd_if_fire_2;
  wire                ll_io_ll_res_if_fire_2;
  wire                when_LockTableBW_l243;
  wire                when_LockTableBW_l252;
  wire                io_lkResp_fire;
  wire                io_lkResp_fire_1;
  `ifndef SYNTHESIS
  reg [47:0] io_lkReq_payload_lkType_string;
  reg [47:0] io_lkResp_payload_lkType_string;
  reg [71:0] io_lkResp_payload_respType_string;
  reg [47:0] htFsm_rLkReq_lkType_string;
  reg [71:0] htFsm_rLkResp_string;
  reg [79:0] htFsm_stateReg_string;
  reg [79:0] htFsm_stateNext_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_string;
  reg [47:0] _zz_htFsm_rLkReq_lkType_1_string;
  reg [47:0] _zz_io_ll_cmd_if_payload_key_string;
  `endif


  assign _zz_htFsm_htNewRamEntry_ownerCnt = (htFsm_htRamEntry_ownerCnt - 8'h01);
  assign _zz_htFsm_htNewRamEntry_ownerCnt_1 = (htFsm_htRamEntry_ownerCnt + 8'h01);
  HashTableBB ht (
    .io_clk_i                         (ht_io_clk_i                              ), //i
    .io_rst_i                         (ht_io_rst_i                              ), //i
    .io_ht_cmd_if_valid               (ht_io_ht_cmd_if_valid                    ), //i
    .io_ht_cmd_if_ready               (ht_io_ht_cmd_if_ready                    ), //o
    .io_ht_cmd_if_payload_key         (ht_io_ht_cmd_if_payload_key[18:0]        ), //i
    .io_ht_cmd_if_payload_value       (ht_io_ht_cmd_if_payload_value[18:0]      ), //i
    .io_ht_cmd_if_payload_opcode      (ht_io_ht_cmd_if_payload_opcode[1:0]      ), //i
    .io_ht_res_if_valid               (ht_io_ht_res_if_valid                    ), //o
    .io_ht_res_if_ready               (1'b1                                     ), //i
    .io_ht_res_if_payload_ram_data    (ht_io_ht_res_if_payload_ram_data[47:0]   ), //o
    .io_ht_res_if_payload_find_addr   (ht_io_ht_res_if_payload_find_addr[8:0]   ), //o
    .io_ht_res_if_payload_chain_state (ht_io_ht_res_if_payload_chain_state[2:0] ), //o
    .io_ht_res_if_payload_found_value (ht_io_ht_res_if_payload_found_value[18:0]), //o
    .io_ht_res_if_payload_bucket      (ht_io_ht_res_if_payload_bucket[7:0]      ), //o
    .io_ht_res_if_payload_rescode     (ht_io_ht_res_if_payload_rescode[2:0]     ), //o
    .io_ht_res_if_payload_opcode      (ht_io_ht_res_if_payload_opcode[1:0]      ), //o
    .io_ht_res_if_payload_value       (ht_io_ht_res_if_payload_value[18:0]      ), //o
    .io_ht_res_if_payload_key         (ht_io_ht_res_if_payload_key[18:0]        ), //o
    .io_ht_clear_ram_run              (1'b0                                     ), //i
    .io_ht_clear_ram_done             (ht_io_ht_clear_ram_done                  ), //o
    .io_dt_clear_ram_run              (1'b0                                     ), //i
    .io_dt_clear_ram_done             (ht_io_dt_clear_ram_done                  ), //o
    .io_update_en                     (ht_io_update_en                          ), //i
    .io_update_data                   (ht_io_update_data[47:0]                  ), //i
    .io_update_addr                   (ht_io_update_addr[8:0]                   ), //i
    .resetn                           (resetn                                   ), //i
    .clk                              (clk                                      )  //i
  );
  LinkedListBB ll (
    .io_clk_i                          (ll_io_clk_i                             ), //i
    .io_rst_i                          (ll_io_rst_i                             ), //i
    .io_ll_cmd_if_valid                (ll_io_ll_cmd_if_valid                   ), //i
    .io_ll_cmd_if_ready                (ll_io_ll_cmd_if_ready                   ), //o
    .io_ll_cmd_if_payload_key          (ll_io_ll_cmd_if_payload_key[43:0]       ), //i
    .io_ll_cmd_if_payload_opcode       (ll_io_ll_cmd_if_payload_opcode[1:0]     ), //i
    .io_ll_cmd_if_payload_head_ptr     (ll_io_ll_cmd_if_payload_head_ptr[8:0]   ), //i
    .io_ll_cmd_if_payload_head_ptr_val (ll_io_ll_cmd_if_payload_head_ptr_val    ), //i
    .io_ll_res_if_valid                (ll_io_ll_res_if_valid                   ), //o
    .io_ll_res_if_ready                (1'b1                                    ), //i
    .io_ll_res_if_payload_key          (ll_io_ll_res_if_payload_key[43:0]       ), //o
    .io_ll_res_if_payload_opcode       (ll_io_ll_res_if_payload_opcode[1:0]     ), //o
    .io_ll_res_if_payload_rescode      (ll_io_ll_res_if_payload_rescode[2:0]    ), //o
    .io_ll_res_if_payload_chain_state  (ll_io_ll_res_if_payload_chain_state[2:0]), //o
    .io_head_table_if_wr_data_ptr      (ll_io_head_table_if_wr_data_ptr[8:0]    ), //o
    .io_head_table_if_wr_data_ptr_val  (ll_io_head_table_if_wr_data_ptr_val     ), //o
    .io_head_table_if_wr_en            (ll_io_head_table_if_wr_en               ), //o
    .io_clear_ram_run_i                (1'b0                                    ), //i
    .io_clear_ram_done_o               (ll_io_clear_ram_done_o                  ), //o
    .resetn                            (resetn                                  ), //i
    .clk                               (clk                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_lkReq_payload_lkType)
      LkT_rd : io_lkReq_payload_lkType_string = "rd    ";
      LkT_wr : io_lkReq_payload_lkType_string = "wr    ";
      LkT_raw : io_lkReq_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkReq_payload_lkType_string = "insTab";
      default : io_lkReq_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_lkType)
      LkT_rd : io_lkResp_payload_lkType_string = "rd    ";
      LkT_wr : io_lkResp_payload_lkType_string = "wr    ";
      LkT_raw : io_lkResp_payload_lkType_string = "raw   ";
      LkT_insTab : io_lkResp_payload_lkType_string = "insTab";
      default : io_lkResp_payload_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_lkResp_payload_respType)
      LockRespType_grant : io_lkResp_payload_respType_string = "grant    ";
      LockRespType_abort : io_lkResp_payload_respType_string = "abort    ";
      LockRespType_waiting : io_lkResp_payload_respType_string = "waiting  ";
      LockRespType_release_1 : io_lkResp_payload_respType_string = "release_1";
      default : io_lkResp_payload_respType_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkReq_lkType)
      LkT_rd : htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : htFsm_rLkReq_lkType_string = "insTab";
      default : htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(htFsm_rLkResp)
      LockRespType_grant : htFsm_rLkResp_string = "grant    ";
      LockRespType_abort : htFsm_rLkResp_string = "abort    ";
      LockRespType_waiting : htFsm_rLkResp_string = "waiting  ";
      LockRespType_release_1 : htFsm_rLkResp_string = "release_1";
      default : htFsm_rLkResp_string = "?????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateReg)
      htFsm_enumDef_BOOT : htFsm_stateReg_string = "BOOT      ";
      htFsm_enumDef_HTINSCMD : htFsm_stateReg_string = "HTINSCMD  ";
      htFsm_enumDef_HTINSRESP : htFsm_stateReg_string = "HTINSRESP ";
      htFsm_enumDef_HTDELCMD : htFsm_stateReg_string = "HTDELCMD  ";
      htFsm_enumDef_HTDELRESP : htFsm_stateReg_string = "HTDELRESP ";
      htFsm_enumDef_LLPUSHCMD : htFsm_stateReg_string = "LLPUSHCMD ";
      htFsm_enumDef_LLPUSHRESP : htFsm_stateReg_string = "LLPUSHRESP";
      htFsm_enumDef_LLPOPCMD : htFsm_stateReg_string = "LLPOPCMD  ";
      htFsm_enumDef_LLPOPRESP : htFsm_stateReg_string = "LLPOPRESP ";
      htFsm_enumDef_LLDELCMD : htFsm_stateReg_string = "LLDELCMD  ";
      htFsm_enumDef_LLDELRESP : htFsm_stateReg_string = "LLDELRESP ";
      htFsm_enumDef_LKRESPPOP : htFsm_stateReg_string = "LKRESPPOP ";
      htFsm_enumDef_LKRESP : htFsm_stateReg_string = "LKRESP    ";
      default : htFsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(htFsm_stateNext)
      htFsm_enumDef_BOOT : htFsm_stateNext_string = "BOOT      ";
      htFsm_enumDef_HTINSCMD : htFsm_stateNext_string = "HTINSCMD  ";
      htFsm_enumDef_HTINSRESP : htFsm_stateNext_string = "HTINSRESP ";
      htFsm_enumDef_HTDELCMD : htFsm_stateNext_string = "HTDELCMD  ";
      htFsm_enumDef_HTDELRESP : htFsm_stateNext_string = "HTDELRESP ";
      htFsm_enumDef_LLPUSHCMD : htFsm_stateNext_string = "LLPUSHCMD ";
      htFsm_enumDef_LLPUSHRESP : htFsm_stateNext_string = "LLPUSHRESP";
      htFsm_enumDef_LLPOPCMD : htFsm_stateNext_string = "LLPOPCMD  ";
      htFsm_enumDef_LLPOPRESP : htFsm_stateNext_string = "LLPOPRESP ";
      htFsm_enumDef_LLDELCMD : htFsm_stateNext_string = "LLDELCMD  ";
      htFsm_enumDef_LLDELRESP : htFsm_stateNext_string = "LLDELRESP ";
      htFsm_enumDef_LKRESPPOP : htFsm_stateNext_string = "LKRESPPOP ";
      htFsm_enumDef_LKRESP : htFsm_stateNext_string = "LKRESP    ";
      default : htFsm_stateNext_string = "??????????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType)
      LkT_rd : _zz_htFsm_rLkReq_lkType_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_htFsm_rLkReq_lkType_1)
      LkT_rd : _zz_htFsm_rLkReq_lkType_1_string = "rd    ";
      LkT_wr : _zz_htFsm_rLkReq_lkType_1_string = "wr    ";
      LkT_raw : _zz_htFsm_rLkReq_lkType_1_string = "raw   ";
      LkT_insTab : _zz_htFsm_rLkReq_lkType_1_string = "insTab";
      default : _zz_htFsm_rLkReq_lkType_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_ll_cmd_if_payload_key)
      LkT_rd : _zz_io_ll_cmd_if_payload_key_string = "rd    ";
      LkT_wr : _zz_io_ll_cmd_if_payload_key_string = "wr    ";
      LkT_raw : _zz_io_ll_cmd_if_payload_key_string = "raw   ";
      LkT_insTab : _zz_io_ll_cmd_if_payload_key_string = "insTab";
      default : _zz_io_ll_cmd_if_payload_key_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    ht_io_ht_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        ht_io_ht_cmd_if_valid = io_lkReq_valid;
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
        ht_io_ht_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_key = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_key = io_lkReq_payload_tId;
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_key = htFsm_rLkReq_tId;
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_value = 19'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_value = {htFsm_tryLkEntry_waitQPtrVld,{htFsm_tryLkEntry_waitQPtr,{htFsm_tryLkEntry_ownerCnt,htFsm_tryLkEntry_lkMode}}};
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_value = 19'h0;
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_ht_cmd_if_payload_opcode = HTOp_sea;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_ins2;
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
        ht_io_ht_cmd_if_payload_opcode = HTOp_del;
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_en = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    ht_io_update_en = 1'b1;
                  end
                end
                HTRet_ins_fail : begin
                end
                default : begin
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                end
                default : begin
                  if(!when_LockTableBW_l140) begin
                    ht_io_update_en = 1'b1;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end
        end
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          ht_io_update_en = ll_io_head_table_if_wr_en;
        end
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            ht_io_update_en = ll_io_head_table_if_wr_en;
          end else begin
            if(!when_LockTableBW_l252) begin
              ht_io_update_en = 1'b1;
            end
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_addr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
        ht_io_update_addr = ht_io_ht_res_if_payload_find_addr;
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        ht_io_update_addr = htFsm_rHtRamAddr;
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ht_io_update_data = 48'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        ht_io_update_data = {htFsm_htNewRamEntry_key,{htFsm_htNewRamEntry_waitQPtrVld,{htFsm_htNewRamEntry_waitQPtr,{htFsm_htNewRamEntry_ownerCnt,{htFsm_htNewRamEntry_lkMode,{htFsm_htNewRamEntry_nextPtr,htFsm_htNewRamEntry_nextPtrVld}}}}}};
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_valid = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
        ll_io_ll_cmd_if_valid = 1'b1;
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_key = 44'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{htFsm_rLkReq_txnAbt,{htFsm_rLkReq_txnTimeOut,{htFsm_rLkReq_lkRelease,{htFsm_rLkReq_lkType,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_key = {htFsm_rLkReq_wLen,{htFsm_rLkReq_lkIdx,{_zz_io_ll_cmd_if_payload_key_3,{_zz_io_ll_cmd_if_payload_key_2,{_zz_io_ll_cmd_if_payload_key_1,{_zz_io_ll_cmd_if_payload_key,{htFsm_rLkReq_txnId,{htFsm_rLkReq_snId,{htFsm_rLkReq_tabId,{htFsm_rLkReq_tId,htFsm_rLkReq_nId}}}}}}}}}};
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_ins;
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_deq;
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_opcode = LLOp_del;
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr = 9'h0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr = htFsm_rHtRamEntry_waitQPtr;
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    ll_io_ll_cmd_if_payload_head_ptr_val = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
        ll_io_ll_cmd_if_payload_head_ptr_val = htFsm_rHtRamEntry_waitQPtrVld;
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_lkReq_ready = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        io_lkReq_ready = ht_io_ht_cmd_if_ready;
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_wantExit = 1'b0;
  always @(*) begin
    htFsm_wantStart = 1'b0;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
        htFsm_wantStart = 1'b1;
      end
    endcase
  end

  assign htFsm_wantKill = 1'b0;
  assign _zz_htFsm_htLkEntry_lkMode = ht_io_ht_res_if_payload_found_value;
  assign htFsm_htLkEntry_lkMode = _zz_htFsm_htLkEntry_lkMode[0];
  assign htFsm_htLkEntry_ownerCnt = _zz_htFsm_htLkEntry_lkMode[8 : 1];
  assign htFsm_htLkEntry_waitQPtr = _zz_htFsm_htLkEntry_lkMode[17 : 9];
  assign htFsm_htLkEntry_waitQPtrVld = _zz_htFsm_htLkEntry_lkMode[18];
  assign _zz_htFsm_htRamEntry_nextPtrVld = ht_io_ht_res_if_payload_ram_data;
  assign htFsm_htRamEntry_nextPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[0];
  assign htFsm_htRamEntry_nextPtr = _zz_htFsm_htRamEntry_nextPtrVld[9 : 1];
  assign htFsm_htRamEntry_lkMode = _zz_htFsm_htRamEntry_nextPtrVld[10];
  assign htFsm_htRamEntry_ownerCnt = _zz_htFsm_htRamEntry_nextPtrVld[18 : 11];
  assign htFsm_htRamEntry_waitQPtr = _zz_htFsm_htRamEntry_nextPtrVld[27 : 19];
  assign htFsm_htRamEntry_waitQPtrVld = _zz_htFsm_htRamEntry_nextPtrVld[28];
  assign htFsm_htRamEntry_key = _zz_htFsm_htRamEntry_nextPtrVld[47 : 29];
  assign ht_io_ht_res_if_fire = (ht_io_ht_res_if_valid && 1'b1);
  assign ht_io_ht_res_if_fire_1 = (ht_io_ht_res_if_valid && 1'b1);
  assign htFsm_htNewRamEntry_nextPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtrVld : htFsm_rHtRamEntry_nextPtrVld);
  assign htFsm_htNewRamEntry_nextPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_nextPtr : htFsm_rHtRamEntry_nextPtr);
  always @(*) begin
    htFsm_htNewRamEntry_lkMode = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_lkMode : htFsm_rHtRamEntry_lkMode);
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        htFsm_htNewRamEntry_lkMode = ((_zz_htFsm_rLkReq_lkType == LkT_wr) || (_zz_htFsm_rLkReq_lkType == LkT_raw));
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_ownerCnt = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_ownerCnt : htFsm_rHtRamEntry_ownerCnt);
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
        htFsm_htNewRamEntry_ownerCnt = (htFsm_rLkReq_lkRelease ? _zz_htFsm_htNewRamEntry_ownerCnt : _zz_htFsm_htNewRamEntry_ownerCnt_1);
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(!when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_ownerCnt = (htFsm_rHtRamEntry_ownerCnt - 8'h01);
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtr = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtr : htFsm_rHtRamEntry_waitQPtr);
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtr = ll_io_head_table_if_wr_data_ptr;
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    htFsm_htNewRamEntry_waitQPtrVld = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_waitQPtrVld : htFsm_rHtRamEntry_waitQPtrVld);
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
      end
      htFsm_enumDef_HTINSRESP : begin
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_htNewRamEntry_waitQPtrVld = ll_io_head_table_if_wr_data_ptr_val;
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  assign htFsm_htNewRamEntry_key = (_zz_htFsm_htNewRamEntry_nextPtrVld ? htFsm_htRamEntry_key : htFsm_rHtRamEntry_key);
  assign io_lkResp_payload_nId = htFsm_rLkReq_nId;
  assign io_lkResp_payload_tId = htFsm_rLkReq_tId;
  assign io_lkResp_payload_tabId = htFsm_rLkReq_tabId;
  assign io_lkResp_payload_snId = htFsm_rLkReq_snId;
  assign io_lkResp_payload_txnId = htFsm_rLkReq_txnId;
  assign io_lkResp_payload_lkType = htFsm_rLkReq_lkType;
  assign io_lkResp_payload_lkRelease = htFsm_rLkReq_lkRelease;
  assign io_lkResp_payload_txnAbt = htFsm_rLkReq_txnAbt;
  assign io_lkResp_payload_lkIdx = htFsm_rLkReq_lkIdx;
  assign io_lkResp_payload_wLen = htFsm_rLkReq_wLen;
  assign io_lkResp_payload_respType = htFsm_rLkResp;
  assign io_lkResp_payload_lkWaited = htFsm_rLkWaited;
  assign io_lkResp_valid = ((htFsm_stateReg == htFsm_enumDef_LKRESP) || (htFsm_stateReg == htFsm_enumDef_LKRESPPOP));
  assign htFsm_tryLkEntry_ownerCnt = 8'h01;
  assign htFsm_tryLkEntry_waitQPtr = 9'h0;
  assign htFsm_tryLkEntry_waitQPtrVld = 1'b0;
  assign htFsm_tryLkEntry_lkMode = ((io_lkReq_payload_lkType == LkT_wr) || (io_lkReq_payload_lkType == LkT_raw));
  always @(*) begin
    htFsm_stateNext = htFsm_stateReg;
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_stateNext = htFsm_enumDef_HTINSRESP;
        end
      end
      htFsm_enumDef_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(when_LockTableBW_l109) begin
                    htFsm_stateNext = htFsm_enumDef_LLPUSHCMD;
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_LKRESP;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_stateNext = htFsm_enumDef_LKRESP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_LKRESP;
                end
              endcase
            end
            default : begin
              case(htFsm_rLkReq_txnTimeOut)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_LLDELCMD;
                end
                default : begin
                  if(when_LockTableBW_l140) begin
                    case(htFsm_htLkEntry_waitQPtrVld)
                      1'b1 : begin
                        htFsm_stateNext = htFsm_enumDef_LKRESPPOP;
                      end
                      default : begin
                        htFsm_stateNext = htFsm_enumDef_HTDELCMD;
                      end
                    endcase
                  end else begin
                    htFsm_stateNext = htFsm_enumDef_LKRESP;
                  end
                end
              endcase
            end
          endcase
        end
      end
      htFsm_enumDef_HTDELCMD : begin
        if(ht_io_ht_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_HTDELRESP;
        end
      end
      htFsm_enumDef_HTDELRESP : begin
        if(ht_io_ht_res_if_fire_3) begin
          htFsm_stateNext = htFsm_enumDef_LKRESP;
        end
      end
      htFsm_enumDef_LLPUSHCMD : begin
        if(ll_io_ll_cmd_if_fire) begin
          htFsm_stateNext = htFsm_enumDef_LLPUSHRESP;
        end
      end
      htFsm_enumDef_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_stateNext = htFsm_enumDef_LKRESP;
          end else begin
            htFsm_stateNext = htFsm_enumDef_LKRESP;
          end
        end
      end
      htFsm_enumDef_LLPOPCMD : begin
        if(ll_io_ll_cmd_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_LLPOPRESP;
        end
      end
      htFsm_enumDef_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_LKRESP;
        end
      end
      htFsm_enumDef_LLDELCMD : begin
        if(ll_io_ll_cmd_if_fire_2) begin
          htFsm_stateNext = htFsm_enumDef_LLDELRESP;
        end
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_stateNext = htFsm_enumDef_LKRESP;
          end else begin
            if(when_LockTableBW_l252) begin
              case(htFsm_htLkEntry_waitQPtrVld)
                1'b1 : begin
                  htFsm_stateNext = htFsm_enumDef_LKRESPPOP;
                end
                default : begin
                  htFsm_stateNext = htFsm_enumDef_HTDELCMD;
                end
              endcase
            end else begin
              htFsm_stateNext = htFsm_enumDef_LKRESP;
            end
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
        if(io_lkResp_fire) begin
          htFsm_stateNext = htFsm_enumDef_LLPOPCMD;
        end
      end
      htFsm_enumDef_LKRESP : begin
        if(io_lkResp_fire_1) begin
          htFsm_stateNext = htFsm_enumDef_HTINSCMD;
        end
      end
      default : begin
      end
    endcase
    if(htFsm_wantStart) begin
      htFsm_stateNext = htFsm_enumDef_HTINSCMD;
    end
    if(htFsm_wantKill) begin
      htFsm_stateNext = htFsm_enumDef_BOOT;
    end
  end

  assign io_lkReq_fire = (io_lkReq_valid && io_lkReq_ready);
  assign ht_io_ht_res_if_fire_2 = (ht_io_ht_res_if_valid && 1'b1);
  assign when_LockTableBW_l109 = (htFsm_htLkEntry_lkMode || ((htFsm_rLkReq_lkType == LkT_wr) || (htFsm_rLkReq_lkType == LkT_raw)));
  assign when_LockTableBW_l140 = (htFsm_htLkEntry_ownerCnt == 8'h01);
  assign ht_io_ht_cmd_if_fire = (ht_io_ht_cmd_if_valid && ht_io_ht_cmd_if_ready);
  assign ht_io_ht_res_if_fire_3 = (ht_io_ht_res_if_valid && 1'b1);
  assign ll_io_ll_cmd_if_fire = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l184 = (ll_io_ll_res_if_payload_rescode == LLRet_ins_success);
  assign ll_io_ll_cmd_if_fire_1 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign _zz_htFsm_rLkReq_nId = ll_io_ll_res_if_payload_key;
  assign _zz_htFsm_rLkReq_lkType_1 = _zz_htFsm_rLkReq_nId[31 : 30];
  assign _zz_htFsm_rLkReq_lkType = _zz_htFsm_rLkReq_lkType_1;
  assign ll_io_ll_res_if_fire_1 = (ll_io_ll_res_if_valid && 1'b1);
  assign _zz_io_ll_cmd_if_payload_key = htFsm_rLkReq_lkType;
  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_1 = htFsm_rLkReq_lkRelease;
    _zz_io_ll_cmd_if_payload_key_1 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_2 = htFsm_rLkReq_txnTimeOut;
    _zz_io_ll_cmd_if_payload_key_2 = 1'b0;
  end

  always @(*) begin
    _zz_io_ll_cmd_if_payload_key_3 = htFsm_rLkReq_txnAbt;
    _zz_io_ll_cmd_if_payload_key_3 = 1'b0;
  end

  assign ll_io_ll_cmd_if_fire_2 = (ll_io_ll_cmd_if_valid && ll_io_ll_cmd_if_ready);
  assign ll_io_ll_res_if_fire_2 = (ll_io_ll_res_if_valid && 1'b1);
  assign when_LockTableBW_l243 = (ll_io_ll_res_if_payload_rescode == LLRet_del_success);
  assign when_LockTableBW_l252 = (htFsm_rHtRamEntry_ownerCnt == 8'h01);
  assign io_lkResp_fire = (io_lkResp_valid && io_lkResp_ready);
  assign io_lkResp_fire_1 = (io_lkResp_valid && io_lkResp_ready);
  assign _zz_htFsm_htNewRamEntry_nextPtrVld = (htFsm_stateReg == htFsm_enumDef_HTINSRESP);
  always @(posedge clk) begin
    if(ht_io_ht_res_if_fire) begin
      htFsm_rHtRamEntry_nextPtrVld <= htFsm_htRamEntry_nextPtrVld;
      htFsm_rHtRamEntry_nextPtr <= htFsm_htRamEntry_nextPtr;
      htFsm_rHtRamEntry_lkMode <= htFsm_htRamEntry_lkMode;
      htFsm_rHtRamEntry_ownerCnt <= htFsm_htRamEntry_ownerCnt;
      htFsm_rHtRamEntry_waitQPtr <= htFsm_htRamEntry_waitQPtr;
      htFsm_rHtRamEntry_waitQPtrVld <= htFsm_htRamEntry_waitQPtrVld;
      htFsm_rHtRamEntry_key <= htFsm_htRamEntry_key;
    end
    if(ht_io_ht_res_if_fire_1) begin
      htFsm_rHtRamAddr <= ht_io_update_addr;
    end
    case(htFsm_stateReg)
      htFsm_enumDef_HTINSCMD : begin
        if(io_lkReq_fire) begin
          htFsm_rLkReq_nId <= io_lkReq_payload_nId;
          htFsm_rLkReq_tId <= io_lkReq_payload_tId;
          htFsm_rLkReq_tabId <= io_lkReq_payload_tabId;
          htFsm_rLkReq_snId <= io_lkReq_payload_snId;
          htFsm_rLkReq_txnId <= io_lkReq_payload_txnId;
          htFsm_rLkReq_lkType <= io_lkReq_payload_lkType;
          htFsm_rLkReq_lkRelease <= io_lkReq_payload_lkRelease;
          htFsm_rLkReq_txnTimeOut <= io_lkReq_payload_txnTimeOut;
          htFsm_rLkReq_txnAbt <= io_lkReq_payload_txnAbt;
          htFsm_rLkReq_lkIdx <= io_lkReq_payload_lkIdx;
          htFsm_rLkReq_wLen <= io_lkReq_payload_wLen;
        end
      end
      htFsm_enumDef_HTINSRESP : begin
        if(ht_io_ht_res_if_fire_2) begin
          htFsm_rLkWaited <= 1'b0;
          case(htFsm_rLkReq_lkRelease)
            1'b0 : begin
              case(ht_io_ht_res_if_payload_rescode)
                HTRet_ins_exist : begin
                  if(!when_LockTableBW_l109) begin
                    htFsm_rLkResp <= LockRespType_grant;
                  end
                end
                HTRet_ins_fail : begin
                  htFsm_rLkResp <= LockRespType_abort;
                end
                default : begin
                  htFsm_rLkResp <= LockRespType_grant;
                end
              endcase
            end
            default : begin
              htFsm_rLkResp <= LockRespType_release_1;
            end
          endcase
        end
      end
      htFsm_enumDef_HTDELCMD : begin
      end
      htFsm_enumDef_HTDELRESP : begin
      end
      htFsm_enumDef_LLPUSHCMD : begin
      end
      htFsm_enumDef_LLPUSHRESP : begin
        if(ll_io_ll_res_if_fire) begin
          if(when_LockTableBW_l184) begin
            htFsm_rLkResp <= LockRespType_waiting;
          end else begin
            htFsm_rLkResp <= LockRespType_abort;
          end
        end
      end
      htFsm_enumDef_LLPOPCMD : begin
      end
      htFsm_enumDef_LLPOPRESP : begin
        if(ll_io_ll_res_if_fire_1) begin
          htFsm_rLkReq_nId <= _zz_htFsm_rLkReq_nId[0 : 0];
          htFsm_rLkReq_tId <= _zz_htFsm_rLkReq_nId[19 : 1];
          htFsm_rLkReq_tabId <= _zz_htFsm_rLkReq_nId[22 : 20];
          htFsm_rLkReq_snId <= _zz_htFsm_rLkReq_nId[23 : 23];
          htFsm_rLkReq_txnId <= _zz_htFsm_rLkReq_nId[29 : 24];
          htFsm_rLkReq_lkType <= _zz_htFsm_rLkReq_lkType;
          htFsm_rLkReq_lkRelease <= _zz_htFsm_rLkReq_nId[32];
          htFsm_rLkReq_txnTimeOut <= _zz_htFsm_rLkReq_nId[33];
          htFsm_rLkReq_txnAbt <= _zz_htFsm_rLkReq_nId[34];
          htFsm_rLkReq_lkIdx <= _zz_htFsm_rLkReq_nId[40 : 35];
          htFsm_rLkReq_wLen <= _zz_htFsm_rLkReq_nId[43 : 41];
          htFsm_rLkResp <= LockRespType_grant;
          htFsm_rLkWaited <= 1'b1;
        end
      end
      htFsm_enumDef_LLDELCMD : begin
      end
      htFsm_enumDef_LLDELRESP : begin
        if(ll_io_ll_res_if_fire_2) begin
          if(when_LockTableBW_l243) begin
            htFsm_rLkResp <= LockRespType_release_1;
            htFsm_rLkWaited <= 1'b1;
          end
        end
      end
      htFsm_enumDef_LKRESPPOP : begin
      end
      htFsm_enumDef_LKRESP : begin
      end
      default : begin
      end
    endcase
  end

  always @(posedge clk) begin
    if(!resetn) begin
      htFsm_stateReg <= htFsm_enumDef_BOOT;
    end else begin
      htFsm_stateReg <= htFsm_stateNext;
    end
  end


endmodule

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

//LinkedListBB replaced by LinkedListBB

//HashTableBB replaced by HashTableBB

module LinkedListBB (
  input               io_clk_i,
  input               io_rst_i,
  input               io_ll_cmd_if_valid,
  output              io_ll_cmd_if_ready,
  input      [43:0]   io_ll_cmd_if_payload_key,
  input      [1:0]    io_ll_cmd_if_payload_opcode,
  input      [8:0]    io_ll_cmd_if_payload_head_ptr,
  input               io_ll_cmd_if_payload_head_ptr_val,
  output              io_ll_res_if_valid,
  input               io_ll_res_if_ready,
  output     [43:0]   io_ll_res_if_payload_key,
  output     [1:0]    io_ll_res_if_payload_opcode,
  output     [2:0]    io_ll_res_if_payload_rescode,
  output     [2:0]    io_ll_res_if_payload_chain_state,
  output     [8:0]    io_head_table_if_wr_data_ptr,
  output              io_head_table_if_wr_data_ptr_val,
  output              io_head_table_if_wr_en,
  input               io_clear_ram_run_i,
  output              io_clear_ram_done_o,
  input               resetn,
  input               clk
);
  localparam LLOp_ins = 2'd0;
  localparam LLOp_del = 2'd1;
  localparam LLOp_deq = 2'd2;
  localparam LLRet_ins_success = 3'd0;
  localparam LLRet_ins_exist = 3'd1;
  localparam LLRet_ins_fail = 3'd2;
  localparam LLRet_del_success = 3'd3;
  localparam LLRet_del_fail = 3'd4;
  localparam LLRet_deq_success = 3'd5;
  localparam LLRet_deq_fail = 3'd6;

  wire                ll_rst_i;
  wire                ll_ll_cmd_if_ready;
  wire                ll_ll_res_if_valid;
  wire       [43:0]   ll_ll_res_if_key;
  wire       [1:0]    ll_ll_res_if_opcode;
  wire       [2:0]    ll_ll_res_if_rescode;
  wire       [2:0]    ll_ll_res_if_chain_state;
  wire       [8:0]    ll_head_table_if_wr_data_ptr;
  wire                ll_head_table_if_wr_data_ptr_val;
  wire                ll_head_table_if_wr_en;
  wire                ll_clear_ram_done_o;
  `ifndef SYNTHESIS
  reg [23:0] io_ll_cmd_if_payload_opcode_string;
  reg [87:0] io_ll_res_if_payload_rescode_string;
  `endif


  linked_list_top ll (
    .clk_i                         (clk                               ), //i
    .rst_i                         (ll_rst_i                          ), //i
    .ll_cmd_if_valid               (io_ll_cmd_if_valid                ), //i
    .ll_cmd_if_ready               (ll_ll_cmd_if_ready                ), //o
    .ll_cmd_if_key                 (io_ll_cmd_if_payload_key[43:0]    ), //i
    .ll_cmd_if_opcode              (io_ll_cmd_if_payload_opcode[1:0]  ), //i
    .ll_cmd_if_head_ptr            (io_ll_cmd_if_payload_head_ptr[8:0]), //i
    .ll_cmd_if_head_ptr_val        (io_ll_cmd_if_payload_head_ptr_val ), //i
    .ll_res_if_valid               (ll_ll_res_if_valid                ), //o
    .ll_res_if_ready               (io_ll_res_if_ready                ), //i
    .ll_res_if_key                 (ll_ll_res_if_key[43:0]            ), //o
    .ll_res_if_opcode              (ll_ll_res_if_opcode[1:0]          ), //o
    .ll_res_if_rescode             (ll_ll_res_if_rescode[2:0]         ), //o
    .ll_res_if_chain_state         (ll_ll_res_if_chain_state[2:0]     ), //o
    .head_table_if_wr_data_ptr     (ll_head_table_if_wr_data_ptr[8:0] ), //o
    .head_table_if_wr_data_ptr_val (ll_head_table_if_wr_data_ptr_val  ), //o
    .head_table_if_wr_en           (ll_head_table_if_wr_en            ), //o
    .clear_ram_run_i               (1'b0                              ), //i
    .clear_ram_done_o              (ll_clear_ram_done_o               )  //o
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ll_cmd_if_payload_opcode)
      LLOp_ins : io_ll_cmd_if_payload_opcode_string = "ins";
      LLOp_del : io_ll_cmd_if_payload_opcode_string = "del";
      LLOp_deq : io_ll_cmd_if_payload_opcode_string = "deq";
      default : io_ll_cmd_if_payload_opcode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_ll_res_if_payload_rescode)
      LLRet_ins_success : io_ll_res_if_payload_rescode_string = "ins_success";
      LLRet_ins_exist : io_ll_res_if_payload_rescode_string = "ins_exist  ";
      LLRet_ins_fail : io_ll_res_if_payload_rescode_string = "ins_fail   ";
      LLRet_del_success : io_ll_res_if_payload_rescode_string = "del_success";
      LLRet_del_fail : io_ll_res_if_payload_rescode_string = "del_fail   ";
      LLRet_deq_success : io_ll_res_if_payload_rescode_string = "deq_success";
      LLRet_deq_fail : io_ll_res_if_payload_rescode_string = "deq_fail   ";
      default : io_ll_res_if_payload_rescode_string = "???????????";
    endcase
  end
  `endif

  assign ll_rst_i = (! resetn);
  assign io_ll_cmd_if_ready = ll_ll_cmd_if_ready;
  assign io_ll_res_if_valid = ll_ll_res_if_valid;
  assign io_ll_res_if_payload_key = ll_ll_res_if_key;
  assign io_ll_res_if_payload_opcode = ll_ll_res_if_opcode;
  assign io_ll_res_if_payload_rescode = ll_ll_res_if_rescode;
  assign io_ll_res_if_payload_chain_state = ll_ll_res_if_chain_state;
  assign io_head_table_if_wr_data_ptr = ll_head_table_if_wr_data_ptr;
  assign io_head_table_if_wr_data_ptr_val = ll_head_table_if_wr_data_ptr_val;
  assign io_head_table_if_wr_en = ll_head_table_if_wr_en;
  assign io_clear_ram_done_o = ll_clear_ram_done_o;

endmodule

module HashTableBB (
  input               io_clk_i,
  input               io_rst_i,
  input               io_ht_cmd_if_valid,
  output              io_ht_cmd_if_ready,
  input      [18:0]   io_ht_cmd_if_payload_key,
  input      [18:0]   io_ht_cmd_if_payload_value,
  input      [1:0]    io_ht_cmd_if_payload_opcode,
  output              io_ht_res_if_valid,
  input               io_ht_res_if_ready,
  output     [47:0]   io_ht_res_if_payload_ram_data,
  output     [8:0]    io_ht_res_if_payload_find_addr,
  output     [2:0]    io_ht_res_if_payload_chain_state,
  output     [18:0]   io_ht_res_if_payload_found_value,
  output     [7:0]    io_ht_res_if_payload_bucket,
  output     [2:0]    io_ht_res_if_payload_rescode,
  output     [1:0]    io_ht_res_if_payload_opcode,
  output     [18:0]   io_ht_res_if_payload_value,
  output     [18:0]   io_ht_res_if_payload_key,
  input               io_ht_clear_ram_run,
  output              io_ht_clear_ram_done,
  input               io_dt_clear_ram_run,
  output              io_dt_clear_ram_done,
  input               io_update_en,
  input      [47:0]   io_update_data,
  input      [8:0]    io_update_addr,
  input               resetn,
  input               clk
);
  localparam HTOp_sea = 2'd0;
  localparam HTOp_ins = 2'd1;
  localparam HTOp_del = 2'd2;
  localparam HTOp_ins2 = 2'd3;
  localparam HTRet_sea_success = 3'd0;
  localparam HTRet_sea_fail = 3'd1;
  localparam HTRet_ins_success = 3'd2;
  localparam HTRet_ins_exist = 3'd3;
  localparam HTRet_ins_fail = 3'd4;
  localparam HTRet_del_success = 3'd5;
  localparam HTRet_del_fail = 3'd6;

  wire                ht_rst_i;
  wire                ht_ht_cmd_if_ready;
  wire                ht_ht_res_if_valid;
  wire       [47:0]   ht_ht_res_if_ram_data;
  wire       [8:0]    ht_ht_res_if_find_addr;
  wire       [2:0]    ht_ht_res_if_chain_state;
  wire       [18:0]   ht_ht_res_if_found_value;
  wire       [7:0]    ht_ht_res_if_bucket;
  wire       [2:0]    ht_ht_res_if_rescode;
  wire       [1:0]    ht_ht_res_if_opcode;
  wire       [18:0]   ht_ht_res_if_value;
  wire       [18:0]   ht_ht_res_if_key;
  wire                ht_ht_clear_ram_done;
  wire                ht_dt_clear_ram_done;
  `ifndef SYNTHESIS
  reg [31:0] io_ht_cmd_if_payload_opcode_string;
  reg [87:0] io_ht_res_if_payload_rescode_string;
  `endif


  hash_table_top ht (
    .clk_i                 (clk                             ), //i
    .rst_i                 (ht_rst_i                        ), //i
    .ht_cmd_if_valid       (io_ht_cmd_if_valid              ), //i
    .ht_cmd_if_ready       (ht_ht_cmd_if_ready              ), //o
    .ht_cmd_if_key         (io_ht_cmd_if_payload_key[18:0]  ), //i
    .ht_cmd_if_value       (io_ht_cmd_if_payload_value[18:0]), //i
    .ht_cmd_if_opcode      (io_ht_cmd_if_payload_opcode[1:0]), //i
    .ht_res_if_valid       (ht_ht_res_if_valid              ), //o
    .ht_res_if_ready       (io_ht_res_if_ready              ), //i
    .ht_res_if_ram_data    (ht_ht_res_if_ram_data[47:0]     ), //o
    .ht_res_if_find_addr   (ht_ht_res_if_find_addr[8:0]     ), //o
    .ht_res_if_chain_state (ht_ht_res_if_chain_state[2:0]   ), //o
    .ht_res_if_found_value (ht_ht_res_if_found_value[18:0]  ), //o
    .ht_res_if_bucket      (ht_ht_res_if_bucket[7:0]        ), //o
    .ht_res_if_rescode     (ht_ht_res_if_rescode[2:0]       ), //o
    .ht_res_if_opcode      (ht_ht_res_if_opcode[1:0]        ), //o
    .ht_res_if_value       (ht_ht_res_if_value[18:0]        ), //o
    .ht_res_if_key         (ht_ht_res_if_key[18:0]          ), //o
    .ht_clear_ram_run      (io_ht_clear_ram_run             ), //i
    .ht_clear_ram_done     (ht_ht_clear_ram_done            ), //o
    .dt_clear_ram_run      (io_dt_clear_ram_run             ), //i
    .dt_clear_ram_done     (ht_dt_clear_ram_done            ), //o
    .update_en             (io_update_en                    ), //i
    .update_data           (io_update_data[47:0]            ), //i
    .update_addr           (io_update_addr[8:0]             )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_ht_cmd_if_payload_opcode)
      HTOp_sea : io_ht_cmd_if_payload_opcode_string = "sea ";
      HTOp_ins : io_ht_cmd_if_payload_opcode_string = "ins ";
      HTOp_del : io_ht_cmd_if_payload_opcode_string = "del ";
      HTOp_ins2 : io_ht_cmd_if_payload_opcode_string = "ins2";
      default : io_ht_cmd_if_payload_opcode_string = "????";
    endcase
  end
  always @(*) begin
    case(io_ht_res_if_payload_rescode)
      HTRet_sea_success : io_ht_res_if_payload_rescode_string = "sea_success";
      HTRet_sea_fail : io_ht_res_if_payload_rescode_string = "sea_fail   ";
      HTRet_ins_success : io_ht_res_if_payload_rescode_string = "ins_success";
      HTRet_ins_exist : io_ht_res_if_payload_rescode_string = "ins_exist  ";
      HTRet_ins_fail : io_ht_res_if_payload_rescode_string = "ins_fail   ";
      HTRet_del_success : io_ht_res_if_payload_rescode_string = "del_success";
      HTRet_del_fail : io_ht_res_if_payload_rescode_string = "del_fail   ";
      default : io_ht_res_if_payload_rescode_string = "???????????";
    endcase
  end
  `endif

  assign ht_rst_i = (! resetn);
  assign io_ht_cmd_if_ready = ht_ht_cmd_if_ready;
  assign io_ht_res_if_valid = ht_ht_res_if_valid;
  assign io_ht_res_if_payload_ram_data = ht_ht_res_if_ram_data;
  assign io_ht_res_if_payload_find_addr = ht_ht_res_if_find_addr;
  assign io_ht_res_if_payload_chain_state = ht_ht_res_if_chain_state;
  assign io_ht_res_if_payload_found_value = ht_ht_res_if_found_value;
  assign io_ht_res_if_payload_bucket = ht_ht_res_if_bucket;
  assign io_ht_res_if_payload_rescode = ht_ht_res_if_rescode;
  assign io_ht_res_if_payload_opcode = ht_ht_res_if_opcode;
  assign io_ht_res_if_payload_value = ht_ht_res_if_value;
  assign io_ht_res_if_payload_key = ht_ht_res_if_key;
  assign io_ht_clear_ram_done = ht_ht_clear_ram_done;
  assign io_dt_clear_ram_done = ht_dt_clear_ram_done;

endmodule
